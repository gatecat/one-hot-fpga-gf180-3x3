// This is the unpowered netlist.
module user_proj_example (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \Inst_eFPGA_top.FrameData[100] ;
 wire \Inst_eFPGA_top.FrameData[101] ;
 wire \Inst_eFPGA_top.FrameData[102] ;
 wire \Inst_eFPGA_top.FrameData[103] ;
 wire \Inst_eFPGA_top.FrameData[104] ;
 wire \Inst_eFPGA_top.FrameData[105] ;
 wire \Inst_eFPGA_top.FrameData[106] ;
 wire \Inst_eFPGA_top.FrameData[107] ;
 wire \Inst_eFPGA_top.FrameData[108] ;
 wire \Inst_eFPGA_top.FrameData[109] ;
 wire \Inst_eFPGA_top.FrameData[110] ;
 wire \Inst_eFPGA_top.FrameData[111] ;
 wire \Inst_eFPGA_top.FrameData[112] ;
 wire \Inst_eFPGA_top.FrameData[113] ;
 wire \Inst_eFPGA_top.FrameData[114] ;
 wire \Inst_eFPGA_top.FrameData[115] ;
 wire \Inst_eFPGA_top.FrameData[116] ;
 wire \Inst_eFPGA_top.FrameData[117] ;
 wire \Inst_eFPGA_top.FrameData[118] ;
 wire \Inst_eFPGA_top.FrameData[119] ;
 wire \Inst_eFPGA_top.FrameData[120] ;
 wire \Inst_eFPGA_top.FrameData[121] ;
 wire \Inst_eFPGA_top.FrameData[122] ;
 wire \Inst_eFPGA_top.FrameData[123] ;
 wire \Inst_eFPGA_top.FrameData[124] ;
 wire \Inst_eFPGA_top.FrameData[125] ;
 wire \Inst_eFPGA_top.FrameData[126] ;
 wire \Inst_eFPGA_top.FrameData[127] ;
 wire \Inst_eFPGA_top.FrameData[32] ;
 wire \Inst_eFPGA_top.FrameData[33] ;
 wire \Inst_eFPGA_top.FrameData[34] ;
 wire \Inst_eFPGA_top.FrameData[35] ;
 wire \Inst_eFPGA_top.FrameData[36] ;
 wire \Inst_eFPGA_top.FrameData[37] ;
 wire \Inst_eFPGA_top.FrameData[38] ;
 wire \Inst_eFPGA_top.FrameData[39] ;
 wire \Inst_eFPGA_top.FrameData[40] ;
 wire \Inst_eFPGA_top.FrameData[41] ;
 wire \Inst_eFPGA_top.FrameData[42] ;
 wire \Inst_eFPGA_top.FrameData[43] ;
 wire \Inst_eFPGA_top.FrameData[44] ;
 wire \Inst_eFPGA_top.FrameData[45] ;
 wire \Inst_eFPGA_top.FrameData[46] ;
 wire \Inst_eFPGA_top.FrameData[47] ;
 wire \Inst_eFPGA_top.FrameData[48] ;
 wire \Inst_eFPGA_top.FrameData[49] ;
 wire \Inst_eFPGA_top.FrameData[50] ;
 wire \Inst_eFPGA_top.FrameData[51] ;
 wire \Inst_eFPGA_top.FrameData[52] ;
 wire \Inst_eFPGA_top.FrameData[53] ;
 wire \Inst_eFPGA_top.FrameData[54] ;
 wire \Inst_eFPGA_top.FrameData[55] ;
 wire \Inst_eFPGA_top.FrameData[56] ;
 wire \Inst_eFPGA_top.FrameData[57] ;
 wire \Inst_eFPGA_top.FrameData[58] ;
 wire \Inst_eFPGA_top.FrameData[59] ;
 wire \Inst_eFPGA_top.FrameData[60] ;
 wire \Inst_eFPGA_top.FrameData[61] ;
 wire \Inst_eFPGA_top.FrameData[62] ;
 wire \Inst_eFPGA_top.FrameData[63] ;
 wire \Inst_eFPGA_top.FrameData[64] ;
 wire \Inst_eFPGA_top.FrameData[65] ;
 wire \Inst_eFPGA_top.FrameData[66] ;
 wire \Inst_eFPGA_top.FrameData[67] ;
 wire \Inst_eFPGA_top.FrameData[68] ;
 wire \Inst_eFPGA_top.FrameData[69] ;
 wire \Inst_eFPGA_top.FrameData[70] ;
 wire \Inst_eFPGA_top.FrameData[71] ;
 wire \Inst_eFPGA_top.FrameData[72] ;
 wire \Inst_eFPGA_top.FrameData[73] ;
 wire \Inst_eFPGA_top.FrameData[74] ;
 wire \Inst_eFPGA_top.FrameData[75] ;
 wire \Inst_eFPGA_top.FrameData[76] ;
 wire \Inst_eFPGA_top.FrameData[77] ;
 wire \Inst_eFPGA_top.FrameData[78] ;
 wire \Inst_eFPGA_top.FrameData[79] ;
 wire \Inst_eFPGA_top.FrameData[80] ;
 wire \Inst_eFPGA_top.FrameData[81] ;
 wire \Inst_eFPGA_top.FrameData[82] ;
 wire \Inst_eFPGA_top.FrameData[83] ;
 wire \Inst_eFPGA_top.FrameData[84] ;
 wire \Inst_eFPGA_top.FrameData[85] ;
 wire \Inst_eFPGA_top.FrameData[86] ;
 wire \Inst_eFPGA_top.FrameData[87] ;
 wire \Inst_eFPGA_top.FrameData[88] ;
 wire \Inst_eFPGA_top.FrameData[89] ;
 wire \Inst_eFPGA_top.FrameData[90] ;
 wire \Inst_eFPGA_top.FrameData[91] ;
 wire \Inst_eFPGA_top.FrameData[92] ;
 wire \Inst_eFPGA_top.FrameData[93] ;
 wire \Inst_eFPGA_top.FrameData[94] ;
 wire \Inst_eFPGA_top.FrameData[95] ;
 wire \Inst_eFPGA_top.FrameData[96] ;
 wire \Inst_eFPGA_top.FrameData[97] ;
 wire \Inst_eFPGA_top.FrameData[98] ;
 wire \Inst_eFPGA_top.FrameData[99] ;
 wire \Inst_eFPGA_top.FrameSelect[0] ;
 wire \Inst_eFPGA_top.FrameSelect[100] ;
 wire \Inst_eFPGA_top.FrameSelect[101] ;
 wire \Inst_eFPGA_top.FrameSelect[102] ;
 wire \Inst_eFPGA_top.FrameSelect[103] ;
 wire \Inst_eFPGA_top.FrameSelect[104] ;
 wire \Inst_eFPGA_top.FrameSelect[105] ;
 wire \Inst_eFPGA_top.FrameSelect[106] ;
 wire \Inst_eFPGA_top.FrameSelect[107] ;
 wire \Inst_eFPGA_top.FrameSelect[108] ;
 wire \Inst_eFPGA_top.FrameSelect[109] ;
 wire \Inst_eFPGA_top.FrameSelect[10] ;
 wire \Inst_eFPGA_top.FrameSelect[110] ;
 wire \Inst_eFPGA_top.FrameSelect[111] ;
 wire \Inst_eFPGA_top.FrameSelect[112] ;
 wire \Inst_eFPGA_top.FrameSelect[113] ;
 wire \Inst_eFPGA_top.FrameSelect[114] ;
 wire \Inst_eFPGA_top.FrameSelect[115] ;
 wire \Inst_eFPGA_top.FrameSelect[116] ;
 wire \Inst_eFPGA_top.FrameSelect[117] ;
 wire \Inst_eFPGA_top.FrameSelect[118] ;
 wire \Inst_eFPGA_top.FrameSelect[119] ;
 wire \Inst_eFPGA_top.FrameSelect[11] ;
 wire \Inst_eFPGA_top.FrameSelect[120] ;
 wire \Inst_eFPGA_top.FrameSelect[121] ;
 wire \Inst_eFPGA_top.FrameSelect[122] ;
 wire \Inst_eFPGA_top.FrameSelect[123] ;
 wire \Inst_eFPGA_top.FrameSelect[124] ;
 wire \Inst_eFPGA_top.FrameSelect[125] ;
 wire \Inst_eFPGA_top.FrameSelect[126] ;
 wire \Inst_eFPGA_top.FrameSelect[127] ;
 wire \Inst_eFPGA_top.FrameSelect[128] ;
 wire \Inst_eFPGA_top.FrameSelect[129] ;
 wire \Inst_eFPGA_top.FrameSelect[12] ;
 wire \Inst_eFPGA_top.FrameSelect[130] ;
 wire \Inst_eFPGA_top.FrameSelect[131] ;
 wire \Inst_eFPGA_top.FrameSelect[132] ;
 wire \Inst_eFPGA_top.FrameSelect[133] ;
 wire \Inst_eFPGA_top.FrameSelect[134] ;
 wire \Inst_eFPGA_top.FrameSelect[135] ;
 wire \Inst_eFPGA_top.FrameSelect[136] ;
 wire \Inst_eFPGA_top.FrameSelect[137] ;
 wire \Inst_eFPGA_top.FrameSelect[138] ;
 wire \Inst_eFPGA_top.FrameSelect[139] ;
 wire \Inst_eFPGA_top.FrameSelect[13] ;
 wire \Inst_eFPGA_top.FrameSelect[140] ;
 wire \Inst_eFPGA_top.FrameSelect[141] ;
 wire \Inst_eFPGA_top.FrameSelect[142] ;
 wire \Inst_eFPGA_top.FrameSelect[143] ;
 wire \Inst_eFPGA_top.FrameSelect[144] ;
 wire \Inst_eFPGA_top.FrameSelect[145] ;
 wire \Inst_eFPGA_top.FrameSelect[146] ;
 wire \Inst_eFPGA_top.FrameSelect[147] ;
 wire \Inst_eFPGA_top.FrameSelect[148] ;
 wire \Inst_eFPGA_top.FrameSelect[149] ;
 wire \Inst_eFPGA_top.FrameSelect[14] ;
 wire \Inst_eFPGA_top.FrameSelect[150] ;
 wire \Inst_eFPGA_top.FrameSelect[151] ;
 wire \Inst_eFPGA_top.FrameSelect[152] ;
 wire \Inst_eFPGA_top.FrameSelect[153] ;
 wire \Inst_eFPGA_top.FrameSelect[154] ;
 wire \Inst_eFPGA_top.FrameSelect[155] ;
 wire \Inst_eFPGA_top.FrameSelect[156] ;
 wire \Inst_eFPGA_top.FrameSelect[157] ;
 wire \Inst_eFPGA_top.FrameSelect[158] ;
 wire \Inst_eFPGA_top.FrameSelect[159] ;
 wire \Inst_eFPGA_top.FrameSelect[15] ;
 wire \Inst_eFPGA_top.FrameSelect[160] ;
 wire \Inst_eFPGA_top.FrameSelect[161] ;
 wire \Inst_eFPGA_top.FrameSelect[162] ;
 wire \Inst_eFPGA_top.FrameSelect[163] ;
 wire \Inst_eFPGA_top.FrameSelect[164] ;
 wire \Inst_eFPGA_top.FrameSelect[165] ;
 wire \Inst_eFPGA_top.FrameSelect[166] ;
 wire \Inst_eFPGA_top.FrameSelect[167] ;
 wire \Inst_eFPGA_top.FrameSelect[168] ;
 wire \Inst_eFPGA_top.FrameSelect[169] ;
 wire \Inst_eFPGA_top.FrameSelect[16] ;
 wire \Inst_eFPGA_top.FrameSelect[170] ;
 wire \Inst_eFPGA_top.FrameSelect[171] ;
 wire \Inst_eFPGA_top.FrameSelect[172] ;
 wire \Inst_eFPGA_top.FrameSelect[173] ;
 wire \Inst_eFPGA_top.FrameSelect[174] ;
 wire \Inst_eFPGA_top.FrameSelect[175] ;
 wire \Inst_eFPGA_top.FrameSelect[176] ;
 wire \Inst_eFPGA_top.FrameSelect[177] ;
 wire \Inst_eFPGA_top.FrameSelect[178] ;
 wire \Inst_eFPGA_top.FrameSelect[179] ;
 wire \Inst_eFPGA_top.FrameSelect[17] ;
 wire \Inst_eFPGA_top.FrameSelect[18] ;
 wire \Inst_eFPGA_top.FrameSelect[19] ;
 wire \Inst_eFPGA_top.FrameSelect[1] ;
 wire \Inst_eFPGA_top.FrameSelect[20] ;
 wire \Inst_eFPGA_top.FrameSelect[21] ;
 wire \Inst_eFPGA_top.FrameSelect[22] ;
 wire \Inst_eFPGA_top.FrameSelect[23] ;
 wire \Inst_eFPGA_top.FrameSelect[24] ;
 wire \Inst_eFPGA_top.FrameSelect[25] ;
 wire \Inst_eFPGA_top.FrameSelect[26] ;
 wire \Inst_eFPGA_top.FrameSelect[27] ;
 wire \Inst_eFPGA_top.FrameSelect[28] ;
 wire \Inst_eFPGA_top.FrameSelect[29] ;
 wire \Inst_eFPGA_top.FrameSelect[2] ;
 wire \Inst_eFPGA_top.FrameSelect[30] ;
 wire \Inst_eFPGA_top.FrameSelect[31] ;
 wire \Inst_eFPGA_top.FrameSelect[32] ;
 wire \Inst_eFPGA_top.FrameSelect[33] ;
 wire \Inst_eFPGA_top.FrameSelect[34] ;
 wire \Inst_eFPGA_top.FrameSelect[35] ;
 wire \Inst_eFPGA_top.FrameSelect[36] ;
 wire \Inst_eFPGA_top.FrameSelect[37] ;
 wire \Inst_eFPGA_top.FrameSelect[38] ;
 wire \Inst_eFPGA_top.FrameSelect[39] ;
 wire \Inst_eFPGA_top.FrameSelect[3] ;
 wire \Inst_eFPGA_top.FrameSelect[40] ;
 wire \Inst_eFPGA_top.FrameSelect[41] ;
 wire \Inst_eFPGA_top.FrameSelect[42] ;
 wire \Inst_eFPGA_top.FrameSelect[43] ;
 wire \Inst_eFPGA_top.FrameSelect[44] ;
 wire \Inst_eFPGA_top.FrameSelect[45] ;
 wire \Inst_eFPGA_top.FrameSelect[46] ;
 wire \Inst_eFPGA_top.FrameSelect[47] ;
 wire \Inst_eFPGA_top.FrameSelect[48] ;
 wire \Inst_eFPGA_top.FrameSelect[49] ;
 wire \Inst_eFPGA_top.FrameSelect[4] ;
 wire \Inst_eFPGA_top.FrameSelect[50] ;
 wire \Inst_eFPGA_top.FrameSelect[51] ;
 wire \Inst_eFPGA_top.FrameSelect[52] ;
 wire \Inst_eFPGA_top.FrameSelect[53] ;
 wire \Inst_eFPGA_top.FrameSelect[54] ;
 wire \Inst_eFPGA_top.FrameSelect[55] ;
 wire \Inst_eFPGA_top.FrameSelect[56] ;
 wire \Inst_eFPGA_top.FrameSelect[57] ;
 wire \Inst_eFPGA_top.FrameSelect[58] ;
 wire \Inst_eFPGA_top.FrameSelect[59] ;
 wire \Inst_eFPGA_top.FrameSelect[5] ;
 wire \Inst_eFPGA_top.FrameSelect[60] ;
 wire \Inst_eFPGA_top.FrameSelect[61] ;
 wire \Inst_eFPGA_top.FrameSelect[62] ;
 wire \Inst_eFPGA_top.FrameSelect[63] ;
 wire \Inst_eFPGA_top.FrameSelect[64] ;
 wire \Inst_eFPGA_top.FrameSelect[65] ;
 wire \Inst_eFPGA_top.FrameSelect[66] ;
 wire \Inst_eFPGA_top.FrameSelect[67] ;
 wire \Inst_eFPGA_top.FrameSelect[68] ;
 wire \Inst_eFPGA_top.FrameSelect[69] ;
 wire \Inst_eFPGA_top.FrameSelect[6] ;
 wire \Inst_eFPGA_top.FrameSelect[70] ;
 wire \Inst_eFPGA_top.FrameSelect[71] ;
 wire \Inst_eFPGA_top.FrameSelect[72] ;
 wire \Inst_eFPGA_top.FrameSelect[73] ;
 wire \Inst_eFPGA_top.FrameSelect[74] ;
 wire \Inst_eFPGA_top.FrameSelect[75] ;
 wire \Inst_eFPGA_top.FrameSelect[76] ;
 wire \Inst_eFPGA_top.FrameSelect[77] ;
 wire \Inst_eFPGA_top.FrameSelect[78] ;
 wire \Inst_eFPGA_top.FrameSelect[79] ;
 wire \Inst_eFPGA_top.FrameSelect[7] ;
 wire \Inst_eFPGA_top.FrameSelect[80] ;
 wire \Inst_eFPGA_top.FrameSelect[81] ;
 wire \Inst_eFPGA_top.FrameSelect[82] ;
 wire \Inst_eFPGA_top.FrameSelect[83] ;
 wire \Inst_eFPGA_top.FrameSelect[84] ;
 wire \Inst_eFPGA_top.FrameSelect[85] ;
 wire \Inst_eFPGA_top.FrameSelect[86] ;
 wire \Inst_eFPGA_top.FrameSelect[87] ;
 wire \Inst_eFPGA_top.FrameSelect[88] ;
 wire \Inst_eFPGA_top.FrameSelect[89] ;
 wire \Inst_eFPGA_top.FrameSelect[8] ;
 wire \Inst_eFPGA_top.FrameSelect[90] ;
 wire \Inst_eFPGA_top.FrameSelect[91] ;
 wire \Inst_eFPGA_top.FrameSelect[92] ;
 wire \Inst_eFPGA_top.FrameSelect[93] ;
 wire \Inst_eFPGA_top.FrameSelect[94] ;
 wire \Inst_eFPGA_top.FrameSelect[95] ;
 wire \Inst_eFPGA_top.FrameSelect[96] ;
 wire \Inst_eFPGA_top.FrameSelect[97] ;
 wire \Inst_eFPGA_top.FrameSelect[98] ;
 wire \Inst_eFPGA_top.FrameSelect[99] ;
 wire \Inst_eFPGA_top.FrameSelect[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_Co ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_I_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_T_top ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_config_C_bit0 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_config_C_bit1 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_config_C_bit2 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_config_C_bit3 ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[16] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[17] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[18] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[19] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[20] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[21] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[22] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[23] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[24] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[25] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[26] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[27] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[28] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[29] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[30] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[31] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[32] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[33] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[34] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[35] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_OutputEnable_O ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_UserCLKo ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[9] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[0] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[10] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[11] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[12] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[13] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[14] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[15] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[1] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[2] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[3] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[4] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[5] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[6] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[7] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[8] ;
 wire \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire \fstb_ctr[0] ;
 wire \fstb_ctr[10] ;
 wire \fstb_ctr[11] ;
 wire \fstb_ctr[12] ;
 wire \fstb_ctr[13] ;
 wire \fstb_ctr[14] ;
 wire \fstb_ctr[15] ;
 wire \fstb_ctr[1] ;
 wire \fstb_ctr[2] ;
 wire \fstb_ctr[3] ;
 wire \fstb_ctr[4] ;
 wire \fstb_ctr[5] ;
 wire \fstb_ctr[6] ;
 wire \fstb_ctr[7] ;
 wire \fstb_ctr[8] ;
 wire \fstb_ctr[9] ;
 wire net186;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net187;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net67;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net68;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net91;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net92;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net93;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net94;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net153;
 wire net154;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net155;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net156;
 wire net184;
 wire net185;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire [5:0] clknet_0_io_in;
 wire [5:0] clknet_2_0_0_io_in;
 wire [5:0] clknet_2_1_0_io_in;
 wire [5:0] clknet_2_2_0_io_in;
 wire [5:0] clknet_2_3_0_io_in;
 wire [5:0] clknet_3_0_0_io_in;
 wire [5:0] clknet_3_0_1_io_in;
 wire [5:0] clknet_3_1_0_io_in;
 wire [5:0] clknet_3_1_1_io_in;
 wire [5:0] clknet_3_2_0_io_in;
 wire [5:0] clknet_3_2_1_io_in;
 wire [5:0] clknet_3_3_0_io_in;
 wire [5:0] clknet_3_3_1_io_in;
 wire [5:0] clknet_3_4_0_io_in;
 wire [5:0] clknet_3_4_1_io_in;
 wire [5:0] clknet_3_5_0_io_in;
 wire [5:0] clknet_3_5_1_io_in;
 wire [5:0] clknet_3_6_0_io_in;
 wire [5:0] clknet_3_6_1_io_in;
 wire [5:0] clknet_3_7_0_io_in;
 wire [5:0] clknet_3_7_1_io_in;
 wire [5:0] clknet_4_0_0_io_in;
 wire [5:0] clknet_4_10_0_io_in;
 wire [5:0] clknet_4_11_0_io_in;
 wire [5:0] clknet_4_12_0_io_in;
 wire [5:0] clknet_4_13_0_io_in;
 wire [5:0] clknet_4_14_0_io_in;
 wire [5:0] clknet_4_15_0_io_in;
 wire [5:0] clknet_4_1_0_io_in;
 wire [5:0] clknet_4_2_0_io_in;
 wire [5:0] clknet_4_3_0_io_in;
 wire [5:0] clknet_4_4_0_io_in;
 wire [5:0] clknet_4_5_0_io_in;
 wire [5:0] clknet_4_6_0_io_in;
 wire [5:0] clknet_4_7_0_io_in;
 wire [5:0] clknet_4_8_0_io_in;
 wire [5:0] clknet_4_9_0_io_in;
 wire [5:0] clknet_opt_1_0_io_in;
 wire [5:0] clknet_opt_1_1_io_in;
 wire [5:0] clknet_opt_1_2_io_in;

 W_IO \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO  (.A_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_I_top ),
    .A_O_top(net17),
    .A_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_T_top ),
    .A_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_config_C_bit0 ),
    .A_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_config_C_bit1 ),
    .A_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_config_C_bit2 ),
    .A_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_config_C_bit3 ),
    .B_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_I_top ),
    .B_O_top(net16),
    .B_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_T_top ),
    .B_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_config_C_bit0 ),
    .B_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_config_C_bit1 ),
    .B_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_config_C_bit2 ),
    .B_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_config_C_bit3 ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.FrameData[63] ,
    \Inst_eFPGA_top.FrameData[62] ,
    \Inst_eFPGA_top.FrameData[61] ,
    \Inst_eFPGA_top.FrameData[60] ,
    \Inst_eFPGA_top.FrameData[59] ,
    \Inst_eFPGA_top.FrameData[58] ,
    \Inst_eFPGA_top.FrameData[57] ,
    \Inst_eFPGA_top.FrameData[56] ,
    \Inst_eFPGA_top.FrameData[55] ,
    \Inst_eFPGA_top.FrameData[54] ,
    \Inst_eFPGA_top.FrameData[53] ,
    \Inst_eFPGA_top.FrameData[52] ,
    \Inst_eFPGA_top.FrameData[51] ,
    \Inst_eFPGA_top.FrameData[50] ,
    \Inst_eFPGA_top.FrameData[49] ,
    \Inst_eFPGA_top.FrameData[48] ,
    \Inst_eFPGA_top.FrameData[47] ,
    \Inst_eFPGA_top.FrameData[46] ,
    \Inst_eFPGA_top.FrameData[45] ,
    \Inst_eFPGA_top.FrameData[44] ,
    \Inst_eFPGA_top.FrameData[43] ,
    \Inst_eFPGA_top.FrameData[42] ,
    \Inst_eFPGA_top.FrameData[41] ,
    \Inst_eFPGA_top.FrameData[40] ,
    \Inst_eFPGA_top.FrameData[39] ,
    \Inst_eFPGA_top.FrameData[38] ,
    \Inst_eFPGA_top.FrameData[37] ,
    \Inst_eFPGA_top.FrameData[36] ,
    \Inst_eFPGA_top.FrameData[35] ,
    \Inst_eFPGA_top.FrameData[34] ,
    \Inst_eFPGA_top.FrameData[33] ,
    \Inst_eFPGA_top.FrameData[32] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameStrobe_O[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[0] }));
 W_IO \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO  (.A_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_I_top ),
    .A_O_top(net13),
    .A_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_T_top ),
    .A_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_config_C_bit0 ),
    .A_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_config_C_bit1 ),
    .A_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_config_C_bit2 ),
    .A_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_config_C_bit3 ),
    .B_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_I_top ),
    .B_O_top(net12),
    .B_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_T_top ),
    .B_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_config_C_bit0 ),
    .B_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_config_C_bit1 ),
    .B_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_config_C_bit2 ),
    .B_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_config_C_bit3 ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.FrameData[95] ,
    \Inst_eFPGA_top.FrameData[94] ,
    \Inst_eFPGA_top.FrameData[93] ,
    \Inst_eFPGA_top.FrameData[92] ,
    \Inst_eFPGA_top.FrameData[91] ,
    \Inst_eFPGA_top.FrameData[90] ,
    \Inst_eFPGA_top.FrameData[89] ,
    \Inst_eFPGA_top.FrameData[88] ,
    \Inst_eFPGA_top.FrameData[87] ,
    \Inst_eFPGA_top.FrameData[86] ,
    \Inst_eFPGA_top.FrameData[85] ,
    \Inst_eFPGA_top.FrameData[84] ,
    \Inst_eFPGA_top.FrameData[83] ,
    \Inst_eFPGA_top.FrameData[82] ,
    \Inst_eFPGA_top.FrameData[81] ,
    \Inst_eFPGA_top.FrameData[80] ,
    \Inst_eFPGA_top.FrameData[79] ,
    \Inst_eFPGA_top.FrameData[78] ,
    \Inst_eFPGA_top.FrameData[77] ,
    \Inst_eFPGA_top.FrameData[76] ,
    \Inst_eFPGA_top.FrameData[75] ,
    \Inst_eFPGA_top.FrameData[74] ,
    \Inst_eFPGA_top.FrameData[73] ,
    \Inst_eFPGA_top.FrameData[72] ,
    \Inst_eFPGA_top.FrameData[71] ,
    \Inst_eFPGA_top.FrameData[70] ,
    \Inst_eFPGA_top.FrameData[69] ,
    \Inst_eFPGA_top.FrameData[68] ,
    \Inst_eFPGA_top.FrameData[67] ,
    \Inst_eFPGA_top.FrameData[66] ,
    \Inst_eFPGA_top.FrameData[65] ,
    \Inst_eFPGA_top.FrameData[64] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameStrobe_O[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[0] }));
 W_IO \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO  (.A_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_I_top ),
    .A_O_top(net9),
    .A_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_T_top ),
    .A_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_config_C_bit0 ),
    .A_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_config_C_bit1 ),
    .A_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_config_C_bit2 ),
    .A_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_config_C_bit3 ),
    .B_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_I_top ),
    .B_O_top(net8),
    .B_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_T_top ),
    .B_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_config_C_bit0 ),
    .B_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_config_C_bit1 ),
    .B_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_config_C_bit2 ),
    .B_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_config_C_bit3 ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_OutputEnable_O ),
    .UserCLK(net50),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.FrameData[127] ,
    \Inst_eFPGA_top.FrameData[126] ,
    \Inst_eFPGA_top.FrameData[125] ,
    \Inst_eFPGA_top.FrameData[124] ,
    \Inst_eFPGA_top.FrameData[123] ,
    \Inst_eFPGA_top.FrameData[122] ,
    \Inst_eFPGA_top.FrameData[121] ,
    \Inst_eFPGA_top.FrameData[120] ,
    \Inst_eFPGA_top.FrameData[119] ,
    \Inst_eFPGA_top.FrameData[118] ,
    \Inst_eFPGA_top.FrameData[117] ,
    \Inst_eFPGA_top.FrameData[116] ,
    \Inst_eFPGA_top.FrameData[115] ,
    \Inst_eFPGA_top.FrameData[114] ,
    \Inst_eFPGA_top.FrameData[113] ,
    \Inst_eFPGA_top.FrameData[112] ,
    \Inst_eFPGA_top.FrameData[111] ,
    \Inst_eFPGA_top.FrameData[110] ,
    \Inst_eFPGA_top.FrameData[109] ,
    \Inst_eFPGA_top.FrameData[108] ,
    \Inst_eFPGA_top.FrameData[107] ,
    \Inst_eFPGA_top.FrameData[106] ,
    \Inst_eFPGA_top.FrameData[105] ,
    \Inst_eFPGA_top.FrameData[104] ,
    \Inst_eFPGA_top.FrameData[103] ,
    \Inst_eFPGA_top.FrameData[102] ,
    \Inst_eFPGA_top.FrameData[101] ,
    \Inst_eFPGA_top.FrameData[100] ,
    \Inst_eFPGA_top.FrameData[99] ,
    \Inst_eFPGA_top.FrameData[98] ,
    \Inst_eFPGA_top.FrameData[97] ,
    \Inst_eFPGA_top.FrameData[96] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.FrameSelect[35] ,
    \Inst_eFPGA_top.FrameSelect[34] ,
    \Inst_eFPGA_top.FrameSelect[33] ,
    \Inst_eFPGA_top.FrameSelect[32] ,
    \Inst_eFPGA_top.FrameSelect[31] ,
    \Inst_eFPGA_top.FrameSelect[30] ,
    \Inst_eFPGA_top.FrameSelect[29] ,
    \Inst_eFPGA_top.FrameSelect[28] ,
    \Inst_eFPGA_top.FrameSelect[27] ,
    \Inst_eFPGA_top.FrameSelect[26] ,
    \Inst_eFPGA_top.FrameSelect[25] ,
    \Inst_eFPGA_top.FrameSelect[24] ,
    \Inst_eFPGA_top.FrameSelect[23] ,
    \Inst_eFPGA_top.FrameSelect[22] ,
    \Inst_eFPGA_top.FrameSelect[21] ,
    \Inst_eFPGA_top.FrameSelect[20] ,
    \Inst_eFPGA_top.FrameSelect[19] ,
    \Inst_eFPGA_top.FrameSelect[18] ,
    \Inst_eFPGA_top.FrameSelect[17] ,
    \Inst_eFPGA_top.FrameSelect[16] ,
    \Inst_eFPGA_top.FrameSelect[15] ,
    \Inst_eFPGA_top.FrameSelect[14] ,
    \Inst_eFPGA_top.FrameSelect[13] ,
    \Inst_eFPGA_top.FrameSelect[12] ,
    \Inst_eFPGA_top.FrameSelect[11] ,
    \Inst_eFPGA_top.FrameSelect[10] ,
    \Inst_eFPGA_top.FrameSelect[9] ,
    \Inst_eFPGA_top.FrameSelect[8] ,
    \Inst_eFPGA_top.FrameSelect[7] ,
    \Inst_eFPGA_top.FrameSelect[6] ,
    \Inst_eFPGA_top.FrameSelect[5] ,
    \Inst_eFPGA_top.FrameSelect[4] ,
    \Inst_eFPGA_top.FrameSelect[3] ,
    \Inst_eFPGA_top.FrameSelect[2] ,
    \Inst_eFPGA_top.FrameSelect[1] ,
    \Inst_eFPGA_top.FrameSelect[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameStrobe_O[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[0] }));
 N_term_single \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_N_term_single  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_Co ),
    .OutputEnable(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_OutputEnable_O ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_UserCLKo ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_UserCLKo ),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_FrameStrobe_O[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[0] }));
 LUT4AB \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_LUT4AB  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_Co ),
    .Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_Co ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[0] }),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E2BEG[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N1BEG[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N2BEGb[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_N4BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_NN4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S2BEG[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y0_SS4BEG[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W1BEG[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W2BEGb[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_W6BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_WW4BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[0] }));
 LUT4AB \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_LUT4AB  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_Co ),
    .Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_Co ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[0] }),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E2BEG[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N1BEG[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N2BEGb[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_N4BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_NN4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S2BEG[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_SS4BEG[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W1BEG[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W2BEGb[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_W6BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_WW4BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[0] }));
 LUT4AB \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_LUT4AB  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_Co ),
    .Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_Co ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[0] }),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E2BEG[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N1BEG[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N2BEGb[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_N4BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_NN4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S2BEG[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_SS4BEG[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W1BEG[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W2BEGb[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_W6BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_WW4BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[0] }));
 S_term_single \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single  (.Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_Co ),
    .OutputEnable(net50),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_OutputEnable_O ),
    .UserCLK(clknet_4_4_0_io_in[5]),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_UserCLKo ),
    .FrameStrobe({\Inst_eFPGA_top.FrameSelect[71] ,
    \Inst_eFPGA_top.FrameSelect[70] ,
    \Inst_eFPGA_top.FrameSelect[69] ,
    \Inst_eFPGA_top.FrameSelect[68] ,
    \Inst_eFPGA_top.FrameSelect[67] ,
    \Inst_eFPGA_top.FrameSelect[66] ,
    \Inst_eFPGA_top.FrameSelect[65] ,
    \Inst_eFPGA_top.FrameSelect[64] ,
    \Inst_eFPGA_top.FrameSelect[63] ,
    \Inst_eFPGA_top.FrameSelect[62] ,
    \Inst_eFPGA_top.FrameSelect[61] ,
    \Inst_eFPGA_top.FrameSelect[60] ,
    \Inst_eFPGA_top.FrameSelect[59] ,
    \Inst_eFPGA_top.FrameSelect[58] ,
    \Inst_eFPGA_top.FrameSelect[57] ,
    \Inst_eFPGA_top.FrameSelect[56] ,
    \Inst_eFPGA_top.FrameSelect[55] ,
    \Inst_eFPGA_top.FrameSelect[54] ,
    \Inst_eFPGA_top.FrameSelect[53] ,
    \Inst_eFPGA_top.FrameSelect[52] ,
    \Inst_eFPGA_top.FrameSelect[51] ,
    \Inst_eFPGA_top.FrameSelect[50] ,
    \Inst_eFPGA_top.FrameSelect[49] ,
    \Inst_eFPGA_top.FrameSelect[48] ,
    \Inst_eFPGA_top.FrameSelect[47] ,
    \Inst_eFPGA_top.FrameSelect[46] ,
    \Inst_eFPGA_top.FrameSelect[45] ,
    \Inst_eFPGA_top.FrameSelect[44] ,
    \Inst_eFPGA_top.FrameSelect[43] ,
    \Inst_eFPGA_top.FrameSelect[42] ,
    \Inst_eFPGA_top.FrameSelect[41] ,
    \Inst_eFPGA_top.FrameSelect[40] ,
    \Inst_eFPGA_top.FrameSelect[39] ,
    \Inst_eFPGA_top.FrameSelect[38] ,
    \Inst_eFPGA_top.FrameSelect[37] ,
    \Inst_eFPGA_top.FrameSelect[36] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N2BEGb[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_NN4BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S1BEG[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S2BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_S4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_SS4BEG[0] }));
 N_term_single \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_N_term_single  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_Co ),
    .OutputEnable(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_OutputEnable_O ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_UserCLKo ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_UserCLKo ),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_FrameStrobe_O[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[0] }));
 LUT4AB \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_LUT4AB  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_Co ),
    .Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_Co ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[0] }),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E2BEG[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y1_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N1BEG[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N2BEGb[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_N4BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_NN4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S2BEG[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y0_SS4BEG[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W1BEG[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W2BEGb[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_W6BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_WW4BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[0] }));
 LUT4AB \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_LUT4AB  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_Co ),
    .Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_Co ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[0] }),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E2BEG[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y2_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N1BEG[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N2BEGb[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_N4BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_NN4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S2BEG[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_SS4BEG[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W1BEG[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W2BEGb[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_W6BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_WW4BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[0] }));
 LUT4AB \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_LUT4AB  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_Co ),
    .Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_Co ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[0] }),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E2BEG[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y3_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N1BEG[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N2BEGb[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_N4BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_NN4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S2BEG[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_SS4BEG[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W1BEG[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W2BEGb[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_W6BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_WW4BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[0] }));
 S_term_single \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single  (.Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_Co ),
    .OutputEnable(net50),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_OutputEnable_O ),
    .UserCLK(clknet_4_6_0_io_in[5]),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_UserCLKo ),
    .FrameStrobe({\Inst_eFPGA_top.FrameSelect[107] ,
    \Inst_eFPGA_top.FrameSelect[106] ,
    \Inst_eFPGA_top.FrameSelect[105] ,
    \Inst_eFPGA_top.FrameSelect[104] ,
    \Inst_eFPGA_top.FrameSelect[103] ,
    \Inst_eFPGA_top.FrameSelect[102] ,
    \Inst_eFPGA_top.FrameSelect[101] ,
    \Inst_eFPGA_top.FrameSelect[100] ,
    \Inst_eFPGA_top.FrameSelect[99] ,
    \Inst_eFPGA_top.FrameSelect[98] ,
    \Inst_eFPGA_top.FrameSelect[97] ,
    \Inst_eFPGA_top.FrameSelect[96] ,
    \Inst_eFPGA_top.FrameSelect[95] ,
    \Inst_eFPGA_top.FrameSelect[94] ,
    \Inst_eFPGA_top.FrameSelect[93] ,
    \Inst_eFPGA_top.FrameSelect[92] ,
    \Inst_eFPGA_top.FrameSelect[91] ,
    \Inst_eFPGA_top.FrameSelect[90] ,
    \Inst_eFPGA_top.FrameSelect[89] ,
    \Inst_eFPGA_top.FrameSelect[88] ,
    \Inst_eFPGA_top.FrameSelect[87] ,
    \Inst_eFPGA_top.FrameSelect[86] ,
    \Inst_eFPGA_top.FrameSelect[85] ,
    \Inst_eFPGA_top.FrameSelect[84] ,
    \Inst_eFPGA_top.FrameSelect[83] ,
    \Inst_eFPGA_top.FrameSelect[82] ,
    \Inst_eFPGA_top.FrameSelect[81] ,
    \Inst_eFPGA_top.FrameSelect[80] ,
    \Inst_eFPGA_top.FrameSelect[79] ,
    \Inst_eFPGA_top.FrameSelect[78] ,
    \Inst_eFPGA_top.FrameSelect[77] ,
    \Inst_eFPGA_top.FrameSelect[76] ,
    \Inst_eFPGA_top.FrameSelect[75] ,
    \Inst_eFPGA_top.FrameSelect[74] ,
    \Inst_eFPGA_top.FrameSelect[73] ,
    \Inst_eFPGA_top.FrameSelect[72] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N2BEGb[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_NN4BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S1BEG[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S2BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_S4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_SS4BEG[0] }));
 N_term_single \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_N_term_single  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_Co ),
    .OutputEnable(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_OutputEnable_O ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_UserCLKo ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_UserCLKo ),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_FrameStrobe_O[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[0] }));
 LUT4AB \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_LUT4AB  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_Co ),
    .Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_Co ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[0] }),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E2BEG[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y1_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N1BEG[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N2BEGb[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_N4BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_NN4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S2BEG[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y0_SS4BEG[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W1BEG[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W2BEGb[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_W6BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_WW4BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[0] }));
 LUT4AB \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_LUT4AB  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_Co ),
    .Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_Co ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[0] }),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E2BEG[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y2_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N1BEG[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N2BEGb[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_N4BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_NN4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S2BEG[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_SS4BEG[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W1BEG[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W2BEGb[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_W6BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_WW4BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[0] }));
 LUT4AB \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_LUT4AB  (.Ci(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_Co ),
    .Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_Co ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_UserCLKo ),
    .E1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[0] }),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E1BEG[0] }),
    .E2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[0] }),
    .E2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E2BEG[0] }),
    .E6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_E6BEG[0] }),
    .EE4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y3_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N1BEG[0] }),
    .N1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N2BEGb[0] }),
    .N2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[0] }),
    .N2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_N4BEG[0] }),
    .N4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_NN4BEG[0] }),
    .NN4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[0] }),
    .S1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S1BEG[0] }),
    .S2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[0] }),
    .S2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S2BEG[0] }),
    .S4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_S4BEG[0] }),
    .SS4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_SS4BEG[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W1BEG[0] }),
    .W1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W2BEGb[0] }),
    .W2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[0] }),
    .W2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_W6BEG[0] }),
    .W6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_WW4BEG[0] }),
    .WW4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[0] }));
 S_term_single \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single  (.Co(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_Co ),
    .OutputEnable(net50),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_OutputEnable_O ),
    .UserCLK(clknet_opt_1_2_io_in[5]),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_UserCLKo ),
    .FrameStrobe({\Inst_eFPGA_top.FrameSelect[143] ,
    \Inst_eFPGA_top.FrameSelect[142] ,
    \Inst_eFPGA_top.FrameSelect[141] ,
    \Inst_eFPGA_top.FrameSelect[140] ,
    \Inst_eFPGA_top.FrameSelect[139] ,
    \Inst_eFPGA_top.FrameSelect[138] ,
    \Inst_eFPGA_top.FrameSelect[137] ,
    \Inst_eFPGA_top.FrameSelect[136] ,
    \Inst_eFPGA_top.FrameSelect[135] ,
    \Inst_eFPGA_top.FrameSelect[134] ,
    \Inst_eFPGA_top.FrameSelect[133] ,
    \Inst_eFPGA_top.FrameSelect[132] ,
    \Inst_eFPGA_top.FrameSelect[131] ,
    \Inst_eFPGA_top.FrameSelect[130] ,
    \Inst_eFPGA_top.FrameSelect[129] ,
    \Inst_eFPGA_top.FrameSelect[128] ,
    \Inst_eFPGA_top.FrameSelect[127] ,
    \Inst_eFPGA_top.FrameSelect[126] ,
    \Inst_eFPGA_top.FrameSelect[125] ,
    \Inst_eFPGA_top.FrameSelect[124] ,
    \Inst_eFPGA_top.FrameSelect[123] ,
    \Inst_eFPGA_top.FrameSelect[122] ,
    \Inst_eFPGA_top.FrameSelect[121] ,
    \Inst_eFPGA_top.FrameSelect[120] ,
    \Inst_eFPGA_top.FrameSelect[119] ,
    \Inst_eFPGA_top.FrameSelect[118] ,
    \Inst_eFPGA_top.FrameSelect[117] ,
    \Inst_eFPGA_top.FrameSelect[116] ,
    \Inst_eFPGA_top.FrameSelect[115] ,
    \Inst_eFPGA_top.FrameSelect[114] ,
    \Inst_eFPGA_top.FrameSelect[113] ,
    \Inst_eFPGA_top.FrameSelect[112] ,
    \Inst_eFPGA_top.FrameSelect[111] ,
    \Inst_eFPGA_top.FrameSelect[110] ,
    \Inst_eFPGA_top.FrameSelect[109] ,
    \Inst_eFPGA_top.FrameSelect[108] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_FrameStrobe_O[0] }),
    .N1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N1BEG[0] }),
    .N2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEG[0] }),
    .N2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N2BEGb[0] }),
    .N4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_N4BEG[0] }),
    .NN4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_NN4BEG[0] }),
    .S1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S1BEG[0] }),
    .S2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEGb[0] }),
    .S2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S2BEG[0] }),
    .S4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_S4BEG[0] }),
    .SS4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_SS4BEG[0] }));
 E_IO \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_E_IO  (.A_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_I_top ),
    .A_O_top(net15),
    .A_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_T_top ),
    .A_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_config_C_bit0 ),
    .A_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_config_C_bit1 ),
    .A_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_config_C_bit2 ),
    .A_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_config_C_bit3 ),
    .B_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_I_top ),
    .B_O_top(net14),
    .B_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_T_top ),
    .B_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_config_C_bit0 ),
    .B_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_config_C_bit1 ),
    .B_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_config_C_bit2 ),
    .B_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_config_C_bit3 ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_UserCLKo ),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E1BEG[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E2BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_E6BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y1_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_FrameStrobe_O[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W2BEGb[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_WW4BEG[0] }));
 E_IO \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_E_IO  (.A_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_I_top ),
    .A_O_top(net11),
    .A_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_T_top ),
    .A_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_config_C_bit0 ),
    .A_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_config_C_bit1 ),
    .A_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_config_C_bit2 ),
    .A_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_config_C_bit3 ),
    .B_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_I_top ),
    .B_O_top(net10),
    .B_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_T_top ),
    .B_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_config_C_bit0 ),
    .B_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_config_C_bit1 ),
    .B_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_config_C_bit2 ),
    .B_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_config_C_bit3 ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_OutputEnable_O ),
    .UserCLK(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_OutputEnable_O ),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_UserCLKo ),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E1BEG[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E2BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_E6BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y2_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[0] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_FrameStrobe_O[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W2BEGb[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_WW4BEG[0] }));
 E_IO \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO  (.A_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_I_top ),
    .A_O_top(net7),
    .A_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_T_top ),
    .A_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_config_C_bit0 ),
    .A_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_config_C_bit1 ),
    .A_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_config_C_bit2 ),
    .A_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_config_C_bit3 ),
    .B_I_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_I_top ),
    .B_O_top(net6),
    .B_T_top(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_T_top ),
    .B_config_C_bit0(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_config_C_bit0 ),
    .B_config_C_bit1(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_config_C_bit1 ),
    .B_config_C_bit2(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_config_C_bit2 ),
    .B_config_C_bit3(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_config_C_bit3 ),
    .OutputEnable_O(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_OutputEnable_O ),
    .UserCLK(net2),
    .UserCLKo(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_UserCLKo ),
    .E1END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E1BEG[0] }),
    .E2END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEGb[0] }),
    .E2MID({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E2BEG[0] }),
    .E6END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_E6BEG[0] }),
    .EE4END({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_EE4BEG[0] }),
    .FrameData({\Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y3_FrameData_O[0] }),
    .FrameData_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameData_O[0] }),
    .FrameStrobe({\Inst_eFPGA_top.FrameSelect[179] ,
    \Inst_eFPGA_top.FrameSelect[178] ,
    \Inst_eFPGA_top.FrameSelect[177] ,
    \Inst_eFPGA_top.FrameSelect[176] ,
    \Inst_eFPGA_top.FrameSelect[175] ,
    \Inst_eFPGA_top.FrameSelect[174] ,
    \Inst_eFPGA_top.FrameSelect[173] ,
    \Inst_eFPGA_top.FrameSelect[172] ,
    \Inst_eFPGA_top.FrameSelect[171] ,
    \Inst_eFPGA_top.FrameSelect[170] ,
    \Inst_eFPGA_top.FrameSelect[169] ,
    \Inst_eFPGA_top.FrameSelect[168] ,
    \Inst_eFPGA_top.FrameSelect[167] ,
    \Inst_eFPGA_top.FrameSelect[166] ,
    \Inst_eFPGA_top.FrameSelect[165] ,
    \Inst_eFPGA_top.FrameSelect[164] ,
    \Inst_eFPGA_top.FrameSelect[163] ,
    \Inst_eFPGA_top.FrameSelect[162] ,
    \Inst_eFPGA_top.FrameSelect[161] ,
    \Inst_eFPGA_top.FrameSelect[160] ,
    \Inst_eFPGA_top.FrameSelect[159] ,
    \Inst_eFPGA_top.FrameSelect[158] ,
    \Inst_eFPGA_top.FrameSelect[157] ,
    \Inst_eFPGA_top.FrameSelect[156] ,
    \Inst_eFPGA_top.FrameSelect[155] ,
    \Inst_eFPGA_top.FrameSelect[154] ,
    \Inst_eFPGA_top.FrameSelect[153] ,
    \Inst_eFPGA_top.FrameSelect[152] ,
    \Inst_eFPGA_top.FrameSelect[151] ,
    \Inst_eFPGA_top.FrameSelect[150] ,
    \Inst_eFPGA_top.FrameSelect[149] ,
    \Inst_eFPGA_top.FrameSelect[148] ,
    \Inst_eFPGA_top.FrameSelect[147] ,
    \Inst_eFPGA_top.FrameSelect[146] ,
    \Inst_eFPGA_top.FrameSelect[145] ,
    \Inst_eFPGA_top.FrameSelect[144] }),
    .FrameStrobe_O({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[35] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[34] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[33] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[32] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[31] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[30] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[29] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[28] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[27] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[26] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[25] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[24] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[23] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[22] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[21] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[20] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[19] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[18] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[17] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[16] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_FrameStrobe_O[0] }),
    .W1BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W1BEG[0] }),
    .W2BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEG[0] }),
    .W2BEGb({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W2BEGb[0] }),
    .W6BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_W6BEG[0] }),
    .WW4BEG({\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[15] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[14] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[13] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[12] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[11] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[10] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[9] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[8] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[7] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[6] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[5] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[4] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[3] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[2] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[1] ,
    \Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_WW4BEG[0] }));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0626_ (.I(\fstb_ctr[5] ),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0627_ (.I(\fstb_ctr[4] ),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0628_ (.I(_0317_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0629_ (.A1(_0316_),
    .A2(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0630_ (.I(\fstb_ctr[7] ),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0631_ (.I(\fstb_ctr[6] ),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0632_ (.A1(_0320_),
    .A2(_0321_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0633_ (.A1(_0319_),
    .A2(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0634_ (.I(_0323_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0635_ (.I(\fstb_ctr[3] ),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0636_ (.I(\fstb_ctr[2] ),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0637_ (.A1(_0325_),
    .A2(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0638_ (.I(\fstb_ctr[1] ),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0639_ (.I(\fstb_ctr[0] ),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _0640_ (.A1(\fstb_ctr[15] ),
    .A2(\fstb_ctr[14] ),
    .A3(\fstb_ctr[11] ),
    .A4(\fstb_ctr[10] ),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _0641_ (.A1(\fstb_ctr[13] ),
    .A2(\fstb_ctr[12] ),
    .A3(\fstb_ctr[9] ),
    .A4(\fstb_ctr[8] ),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0642_ (.A1(_0328_),
    .A2(_0329_),
    .A3(_0330_),
    .A4(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0643_ (.A1(_0327_),
    .A2(_0332_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0644_ (.I(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0645_ (.A1(_0324_),
    .A2(_0334_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0646_ (.I(\fstb_ctr[0] ),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0647_ (.I(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0648_ (.A1(_0328_),
    .A2(_0336_),
    .A3(_0330_),
    .A4(_0331_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0649_ (.A1(_0327_),
    .A2(_0337_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0650_ (.I(_0338_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0651_ (.A1(_0324_),
    .A2(_0339_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0652_ (.I(\fstb_ctr[1] ),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0653_ (.A1(_0340_),
    .A2(_0335_),
    .A3(_0330_),
    .A4(_0331_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0654_ (.A1(_0327_),
    .A2(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0655_ (.I(_0342_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0656_ (.A1(_0324_),
    .A2(_0343_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0657_ (.A1(_0340_),
    .A2(_0336_),
    .A3(_0330_),
    .A4(_0331_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0658_ (.A1(_0327_),
    .A2(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0659_ (.I(_0345_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0660_ (.A1(_0324_),
    .A2(_0346_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0661_ (.I(_0323_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0662_ (.I(_0326_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0663_ (.A1(_0325_),
    .A2(_0348_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0664_ (.A1(_0332_),
    .A2(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0665_ (.I(_0350_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0666_ (.A1(_0347_),
    .A2(_0351_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0667_ (.A1(_0337_),
    .A2(_0349_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0668_ (.I(_0352_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0669_ (.A1(_0347_),
    .A2(_0353_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0670_ (.A1(_0341_),
    .A2(_0349_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0671_ (.I(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0672_ (.A1(_0347_),
    .A2(_0355_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0673_ (.A1(_0344_),
    .A2(_0349_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0674_ (.I(_0356_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0675_ (.A1(_0347_),
    .A2(_0357_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0676_ (.I(_0323_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0677_ (.A1(_0325_),
    .A2(_0348_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0678_ (.A1(_0332_),
    .A2(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0679_ (.I(_0360_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0680_ (.A1(_0358_),
    .A2(_0361_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0681_ (.A1(_0337_),
    .A2(_0359_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0682_ (.I(_0362_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0683_ (.A1(_0358_),
    .A2(_0363_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0684_ (.A1(_0341_),
    .A2(_0359_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0685_ (.I(_0364_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0686_ (.A1(_0358_),
    .A2(_0365_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0687_ (.A1(_0344_),
    .A2(_0359_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0688_ (.I(_0366_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0689_ (.A1(_0358_),
    .A2(_0367_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0690_ (.I(_0323_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0691_ (.A1(\fstb_ctr[3] ),
    .A2(\fstb_ctr[2] ),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0692_ (.I(_0369_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0693_ (.A1(_0332_),
    .A2(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0694_ (.I(_0371_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0695_ (.A1(_0368_),
    .A2(_0372_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0696_ (.A1(_0337_),
    .A2(_0370_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0697_ (.I(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0698_ (.A1(_0368_),
    .A2(_0374_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0699_ (.A1(_0341_),
    .A2(_0370_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0700_ (.I(_0375_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0701_ (.A1(_0368_),
    .A2(_0376_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0702_ (.A1(_0344_),
    .A2(_0370_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0703_ (.I(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0704_ (.A1(_0368_),
    .A2(_0378_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0705_ (.I(_0316_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0706_ (.I(_0317_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0707_ (.A1(_0379_),
    .A2(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0708_ (.A1(_0322_),
    .A2(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0709_ (.I(_0382_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0710_ (.A1(_0334_),
    .A2(_0383_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0711_ (.A1(_0339_),
    .A2(_0383_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0712_ (.A1(_0343_),
    .A2(_0383_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0713_ (.A1(_0346_),
    .A2(_0383_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0714_ (.I(_0382_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0715_ (.A1(_0351_),
    .A2(_0384_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0716_ (.A1(_0353_),
    .A2(_0384_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0717_ (.A1(_0355_),
    .A2(_0384_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0718_ (.A1(_0357_),
    .A2(_0384_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0719_ (.I(_0382_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0720_ (.A1(_0361_),
    .A2(_0385_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0721_ (.A1(_0363_),
    .A2(_0385_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0722_ (.A1(_0365_),
    .A2(_0385_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0723_ (.A1(_0367_),
    .A2(_0385_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0724_ (.I(_0382_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0725_ (.A1(_0372_),
    .A2(_0386_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0726_ (.A1(_0374_),
    .A2(_0386_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0727_ (.A1(_0376_),
    .A2(_0386_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0728_ (.A1(_0378_),
    .A2(_0386_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0729_ (.I(_0316_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0730_ (.A1(_0387_),
    .A2(_0380_),
    .A3(_0322_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0731_ (.I(_0388_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0732_ (.A1(_0334_),
    .A2(_0389_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0733_ (.A1(_0339_),
    .A2(_0389_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0734_ (.A1(_0343_),
    .A2(_0389_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0735_ (.A1(_0346_),
    .A2(_0389_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0736_ (.I(_0388_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0737_ (.A1(_0351_),
    .A2(_0390_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0738_ (.A1(_0353_),
    .A2(_0390_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0739_ (.A1(_0355_),
    .A2(_0390_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0740_ (.A1(_0357_),
    .A2(_0390_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0741_ (.I(_0388_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0742_ (.A1(_0361_),
    .A2(_0391_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0743_ (.A1(_0363_),
    .A2(_0391_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0744_ (.A1(_0365_),
    .A2(_0391_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0745_ (.A1(_0367_),
    .A2(_0391_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0746_ (.I(_0388_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0747_ (.A1(_0372_),
    .A2(_0392_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0748_ (.A1(_0374_),
    .A2(_0392_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0749_ (.A1(_0376_),
    .A2(_0392_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0750_ (.A1(_0378_),
    .A2(_0392_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0751_ (.I(_0321_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0752_ (.A1(_0320_),
    .A2(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0753_ (.A1(_0316_),
    .A2(_0380_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0754_ (.A1(_0394_),
    .A2(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0755_ (.I(_0396_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0756_ (.A1(_0334_),
    .A2(_0397_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0757_ (.A1(_0339_),
    .A2(_0397_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0758_ (.A1(_0343_),
    .A2(_0397_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0759_ (.A1(_0346_),
    .A2(_0397_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0760_ (.I(_0396_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0761_ (.A1(_0351_),
    .A2(_0398_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0762_ (.A1(_0353_),
    .A2(_0398_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0763_ (.A1(_0355_),
    .A2(_0398_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0764_ (.A1(_0357_),
    .A2(_0398_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0765_ (.I(_0396_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0766_ (.A1(_0361_),
    .A2(_0399_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0767_ (.A1(_0363_),
    .A2(_0399_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0768_ (.A1(_0365_),
    .A2(_0399_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0769_ (.A1(_0367_),
    .A2(_0399_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0770_ (.I(_0396_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0771_ (.A1(_0372_),
    .A2(_0400_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0772_ (.A1(_0374_),
    .A2(_0400_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0773_ (.A1(_0376_),
    .A2(_0400_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0774_ (.A1(_0378_),
    .A2(_0400_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0775_ (.I(_0333_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0776_ (.A1(_0322_),
    .A2(_0395_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0777_ (.I(_0402_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0778_ (.A1(_0401_),
    .A2(_0403_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0779_ (.A1(_0319_),
    .A2(_0394_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0780_ (.I(_0404_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0781_ (.A1(_0401_),
    .A2(_0405_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0782_ (.I(_0338_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0783_ (.A1(_0406_),
    .A2(_0405_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0784_ (.I(_0342_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0785_ (.A1(_0407_),
    .A2(_0405_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0786_ (.I(_0345_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0787_ (.A1(_0408_),
    .A2(_0405_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0788_ (.I(_0350_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0789_ (.I(_0409_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0790_ (.I(_0404_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0791_ (.A1(_0410_),
    .A2(_0411_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0792_ (.I(_0352_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0793_ (.I(_0412_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0794_ (.A1(_0413_),
    .A2(_0411_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0795_ (.I(_0354_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0796_ (.I(_0414_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0797_ (.A1(_0415_),
    .A2(_0411_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0798_ (.I(_0356_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0799_ (.I(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0800_ (.A1(_0417_),
    .A2(_0411_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0801_ (.I(_0360_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0802_ (.I(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0803_ (.I(_0404_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0804_ (.A1(_0419_),
    .A2(_0420_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0805_ (.I(_0362_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0806_ (.I(_0421_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0807_ (.A1(_0422_),
    .A2(_0420_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0808_ (.A1(_0406_),
    .A2(_0403_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0809_ (.I(_0364_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0810_ (.I(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0811_ (.A1(_0424_),
    .A2(_0420_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0812_ (.I(_0366_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0813_ (.I(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0814_ (.A1(_0426_),
    .A2(_0420_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0815_ (.I(_0371_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0816_ (.I(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0817_ (.I(_0404_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0818_ (.A1(_0428_),
    .A2(_0429_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0819_ (.I(_0373_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0820_ (.I(_0430_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0821_ (.A1(_0431_),
    .A2(_0429_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0822_ (.I(_0375_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0823_ (.I(_0432_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0824_ (.A1(_0433_),
    .A2(_0429_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0825_ (.I(_0377_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0826_ (.I(_0434_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0827_ (.A1(_0435_),
    .A2(_0429_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0828_ (.A1(_0381_),
    .A2(_0394_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0829_ (.I(_0436_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0830_ (.A1(_0401_),
    .A2(_0437_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0831_ (.A1(_0406_),
    .A2(_0437_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0832_ (.A1(_0407_),
    .A2(_0437_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0833_ (.A1(_0408_),
    .A2(_0437_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0834_ (.A1(_0407_),
    .A2(_0403_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0835_ (.I(_0436_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0836_ (.A1(_0410_),
    .A2(_0438_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0837_ (.A1(_0413_),
    .A2(_0438_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0838_ (.A1(_0415_),
    .A2(_0438_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0839_ (.A1(_0417_),
    .A2(_0438_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0840_ (.I(_0436_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0841_ (.A1(_0419_),
    .A2(_0439_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0842_ (.A1(_0422_),
    .A2(_0439_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0843_ (.A1(_0424_),
    .A2(_0439_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0844_ (.A1(_0426_),
    .A2(_0439_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0845_ (.I(_0436_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0846_ (.A1(_0428_),
    .A2(_0440_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0847_ (.A1(_0431_),
    .A2(_0440_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0848_ (.A1(_0408_),
    .A2(_0403_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0849_ (.A1(_0433_),
    .A2(_0440_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0850_ (.A1(_0435_),
    .A2(_0440_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0851_ (.A1(_0387_),
    .A2(_0380_),
    .A3(_0394_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0852_ (.I(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0853_ (.A1(_0401_),
    .A2(_0442_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0854_ (.A1(_0406_),
    .A2(_0442_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0855_ (.A1(_0407_),
    .A2(_0442_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0856_ (.A1(_0408_),
    .A2(_0442_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0857_ (.I(_0441_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0858_ (.A1(_0410_),
    .A2(_0443_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0859_ (.A1(_0413_),
    .A2(_0443_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0860_ (.A1(_0415_),
    .A2(_0443_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0861_ (.A1(_0417_),
    .A2(_0443_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0862_ (.I(_0402_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0863_ (.A1(_0410_),
    .A2(_0444_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0864_ (.I(_0441_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0865_ (.A1(_0419_),
    .A2(_0445_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0866_ (.A1(_0422_),
    .A2(_0445_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0867_ (.A1(_0424_),
    .A2(_0445_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0868_ (.A1(_0426_),
    .A2(_0445_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0869_ (.I(_0441_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0870_ (.A1(_0428_),
    .A2(_0446_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0871_ (.A1(_0431_),
    .A2(_0446_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0872_ (.A1(_0433_),
    .A2(_0446_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0873_ (.A1(_0435_),
    .A2(_0446_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0874_ (.I(_0333_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0875_ (.A1(_0320_),
    .A2(_0393_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0876_ (.A1(_0395_),
    .A2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0877_ (.I(_0449_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0878_ (.A1(_0447_),
    .A2(_0450_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0879_ (.I(_0338_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0880_ (.A1(_0451_),
    .A2(_0450_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0881_ (.A1(_0413_),
    .A2(_0444_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0882_ (.I(_0342_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0883_ (.A1(_0452_),
    .A2(_0450_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0884_ (.I(_0345_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0885_ (.A1(_0453_),
    .A2(_0450_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0886_ (.I(_0449_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0887_ (.A1(_0409_),
    .A2(_0454_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0888_ (.A1(_0412_),
    .A2(_0454_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0889_ (.A1(_0415_),
    .A2(_0454_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0890_ (.A1(_0417_),
    .A2(_0454_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0891_ (.I(_0449_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0892_ (.A1(_0419_),
    .A2(_0455_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0893_ (.A1(_0422_),
    .A2(_0455_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0894_ (.A1(_0424_),
    .A2(_0455_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0895_ (.A1(_0426_),
    .A2(_0455_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0896_ (.A1(_0414_),
    .A2(_0444_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0897_ (.I(_0449_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0898_ (.A1(_0428_),
    .A2(_0456_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0899_ (.A1(_0431_),
    .A2(_0456_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0900_ (.A1(_0433_),
    .A2(_0456_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0901_ (.A1(_0435_),
    .A2(_0456_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0902_ (.A1(_0319_),
    .A2(_0448_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0903_ (.I(_0457_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0904_ (.A1(_0447_),
    .A2(_0458_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0905_ (.A1(_0451_),
    .A2(_0458_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0906_ (.A1(_0452_),
    .A2(_0458_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0907_ (.A1(_0453_),
    .A2(_0458_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0908_ (.I(_0457_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0909_ (.A1(_0409_),
    .A2(_0459_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0910_ (.A1(_0412_),
    .A2(_0459_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0911_ (.A1(_0416_),
    .A2(_0444_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0912_ (.A1(_0414_),
    .A2(_0459_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0913_ (.A1(_0416_),
    .A2(_0459_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0914_ (.I(_0457_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0915_ (.A1(_0418_),
    .A2(_0460_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0916_ (.A1(_0421_),
    .A2(_0460_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0917_ (.A1(_0423_),
    .A2(_0460_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0918_ (.A1(_0425_),
    .A2(_0460_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0919_ (.I(_0457_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0920_ (.A1(_0427_),
    .A2(_0461_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0921_ (.A1(_0430_),
    .A2(_0461_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0922_ (.A1(_0432_),
    .A2(_0461_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0923_ (.A1(_0434_),
    .A2(_0461_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0924_ (.I(_0402_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0925_ (.A1(_0418_),
    .A2(_0462_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0926_ (.A1(_0381_),
    .A2(_0448_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0927_ (.I(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0928_ (.A1(_0447_),
    .A2(_0464_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0929_ (.A1(_0451_),
    .A2(_0464_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0930_ (.A1(_0452_),
    .A2(_0464_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0931_ (.A1(_0453_),
    .A2(_0464_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0932_ (.I(_0463_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0933_ (.A1(_0409_),
    .A2(_0465_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0934_ (.A1(_0412_),
    .A2(_0465_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0935_ (.A1(_0414_),
    .A2(_0465_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0936_ (.A1(_0416_),
    .A2(_0465_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0937_ (.I(_0463_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0938_ (.A1(_0418_),
    .A2(_0466_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0939_ (.A1(_0421_),
    .A2(_0466_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0940_ (.A1(_0421_),
    .A2(_0462_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0941_ (.A1(_0423_),
    .A2(_0466_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0942_ (.A1(_0425_),
    .A2(_0466_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0943_ (.I(_0463_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0944_ (.A1(_0427_),
    .A2(_0467_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0945_ (.A1(_0430_),
    .A2(_0467_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0946_ (.A1(_0432_),
    .A2(_0467_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0947_ (.A1(_0434_),
    .A2(_0467_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0948_ (.I(\fstb_ctr[4] ),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0949_ (.A1(_0387_),
    .A2(_0468_),
    .A3(_0448_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0950_ (.A1(_0447_),
    .A2(_0469_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0951_ (.A1(_0451_),
    .A2(_0469_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0952_ (.A1(_0452_),
    .A2(_0469_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0953_ (.A1(_0453_),
    .A2(_0469_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0954_ (.A1(_0423_),
    .A2(_0462_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0955_ (.A1(_0425_),
    .A2(_0462_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0956_ (.I(_0402_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0957_ (.A1(_0427_),
    .A2(_0470_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0958_ (.A1(_0430_),
    .A2(_0470_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0959_ (.A1(_0432_),
    .A2(_0470_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0960_ (.A1(_0434_),
    .A2(_0470_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0961_ (.I(net4),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0962_ (.I(net5),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0963_ (.I(net21),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0964_ (.I(net20),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0965_ (.I(_0472_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0966_ (.A1(_0471_),
    .A2(_0329_),
    .B(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0967_ (.A1(_0471_),
    .A2(_0329_),
    .B(_0474_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0968_ (.I(net20),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0969_ (.A1(_0471_),
    .A2(_0329_),
    .B(_0328_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0970_ (.A1(_0471_),
    .A2(_0328_),
    .A3(_0335_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0971_ (.A1(_0475_),
    .A2(_0476_),
    .A3(_0477_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0972_ (.A1(net21),
    .A2(\fstb_ctr[1] ),
    .A3(_0335_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0973_ (.I(_0478_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0974_ (.A1(_0348_),
    .A2(_0479_),
    .B(_0473_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0975_ (.A1(_0348_),
    .A2(_0479_),
    .B(_0480_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0976_ (.I(net20),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0977_ (.A1(_0326_),
    .A2(_0477_),
    .B(_0325_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0978_ (.A1(\fstb_ctr[3] ),
    .A2(_0326_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0979_ (.A1(_0483_),
    .A2(_0479_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0980_ (.A1(_0481_),
    .A2(_0482_),
    .A3(_0484_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0981_ (.A1(_0468_),
    .A2(_0484_),
    .B(_0473_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0982_ (.A1(_0468_),
    .A2(_0484_),
    .B(_0485_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0983_ (.A1(_0468_),
    .A2(_0484_),
    .B(_0387_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0984_ (.A1(_0379_),
    .A2(_0318_),
    .A3(_0483_),
    .A4(_0478_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0985_ (.A1(_0481_),
    .A2(_0486_),
    .A3(_0487_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0986_ (.A1(_0393_),
    .A2(_0487_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0987_ (.A1(_0475_),
    .A2(_0488_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0988_ (.A1(_0321_),
    .A2(_0487_),
    .B(_0320_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0989_ (.A1(\fstb_ctr[7] ),
    .A2(_0321_),
    .A3(\fstb_ctr[5] ),
    .A4(_0317_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0990_ (.A1(_0483_),
    .A2(_0478_),
    .A3(_0490_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0991_ (.A1(_0481_),
    .A2(_0489_),
    .A3(_0491_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0992_ (.I(\fstb_ctr[8] ),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0993_ (.A1(_0492_),
    .A2(_0491_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0994_ (.A1(_0475_),
    .A2(_0493_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0995_ (.I(\fstb_ctr[9] ),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0996_ (.A1(_0494_),
    .A2(_0492_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0997_ (.A1(_0483_),
    .A2(_0479_),
    .A3(_0490_),
    .A4(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0998_ (.A1(_0494_),
    .A2(_0492_),
    .B(_0472_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0999_ (.A1(_0494_),
    .A2(_0491_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1000_ (.A1(_0496_),
    .A2(_0497_),
    .A3(_0498_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1001_ (.I(\fstb_ctr[10] ),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1002_ (.A1(_0499_),
    .A2(_0496_),
    .B(_0472_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1003_ (.A1(_0499_),
    .A2(_0496_),
    .B(_0500_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1004_ (.A1(_0499_),
    .A2(_0496_),
    .B(\fstb_ctr[11] ),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1005_ (.A1(\fstb_ctr[7] ),
    .A2(\fstb_ctr[6] ),
    .A3(\fstb_ctr[5] ),
    .A4(_0317_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1006_ (.A1(\fstb_ctr[11] ),
    .A2(_0499_),
    .A3(_0494_),
    .A4(_0492_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1007_ (.A1(_0369_),
    .A2(_0477_),
    .A3(_0502_),
    .A4(_0503_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1008_ (.I(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1009_ (.A1(_0481_),
    .A2(_0501_),
    .A3(_0505_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1010_ (.I(\fstb_ctr[12] ),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1011_ (.A1(_0369_),
    .A2(_0477_),
    .A3(_0502_),
    .A4(_0503_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1012_ (.A1(_0506_),
    .A2(_0507_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1013_ (.A1(_0475_),
    .A2(_0508_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1014_ (.I(\fstb_ctr[13] ),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1015_ (.A1(_0509_),
    .A2(_0506_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1016_ (.A1(_0509_),
    .A2(_0506_),
    .B(_0472_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1017_ (.A1(_0509_),
    .A2(_0505_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1018_ (.A1(_0505_),
    .A2(_0510_),
    .B(_0511_),
    .C(_0512_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1019_ (.A1(_0505_),
    .A2(_0510_),
    .B(\fstb_ctr[14] ),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1020_ (.I(\fstb_ctr[14] ),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1021_ (.A1(_0509_),
    .A2(_0506_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1022_ (.A1(_0514_),
    .A2(_0507_),
    .A3(_0515_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1023_ (.A1(net20),
    .A2(_0513_),
    .A3(_0516_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1024_ (.I(\fstb_ctr[15] ),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1025_ (.A1(_0514_),
    .A2(_0507_),
    .A3(_0515_),
    .B(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1026_ (.A1(\fstb_ctr[15] ),
    .A2(\fstb_ctr[14] ),
    .A3(_0504_),
    .A4(_0510_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1027_ (.A1(_0473_),
    .A2(_0518_),
    .A3(_0519_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1028_ (.I(_0520_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1029_ (.I(net18),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1030_ (.I(_0521_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1031_ (.I(_0522_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1032_ (.I0(\Inst_eFPGA_top.FrameData[32] ),
    .I1(\Inst_eFPGA_top.FrameData[33] ),
    .S(_0523_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1033_ (.I(_0524_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1034_ (.I0(\Inst_eFPGA_top.FrameData[33] ),
    .I1(\Inst_eFPGA_top.FrameData[34] ),
    .S(_0523_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1035_ (.I(_0525_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1036_ (.I0(\Inst_eFPGA_top.FrameData[34] ),
    .I1(\Inst_eFPGA_top.FrameData[35] ),
    .S(_0523_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1037_ (.I(_0526_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1038_ (.I0(\Inst_eFPGA_top.FrameData[35] ),
    .I1(\Inst_eFPGA_top.FrameData[36] ),
    .S(_0523_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1039_ (.I(_0527_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1040_ (.I(_0522_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1041_ (.I0(\Inst_eFPGA_top.FrameData[36] ),
    .I1(\Inst_eFPGA_top.FrameData[37] ),
    .S(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1042_ (.I(_0529_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1043_ (.I0(\Inst_eFPGA_top.FrameData[37] ),
    .I1(\Inst_eFPGA_top.FrameData[38] ),
    .S(_0528_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1044_ (.I(_0530_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1045_ (.I0(\Inst_eFPGA_top.FrameData[38] ),
    .I1(\Inst_eFPGA_top.FrameData[39] ),
    .S(_0528_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1046_ (.I(_0531_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1047_ (.I0(\Inst_eFPGA_top.FrameData[39] ),
    .I1(\Inst_eFPGA_top.FrameData[40] ),
    .S(_0528_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1048_ (.I(_0532_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1049_ (.I(_0522_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1050_ (.I0(\Inst_eFPGA_top.FrameData[40] ),
    .I1(\Inst_eFPGA_top.FrameData[41] ),
    .S(_0533_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1051_ (.I(_0534_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1052_ (.I0(\Inst_eFPGA_top.FrameData[41] ),
    .I1(\Inst_eFPGA_top.FrameData[42] ),
    .S(_0533_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1053_ (.I(_0535_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1054_ (.I0(\Inst_eFPGA_top.FrameData[42] ),
    .I1(\Inst_eFPGA_top.FrameData[43] ),
    .S(_0533_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1055_ (.I(_0536_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1056_ (.I0(\Inst_eFPGA_top.FrameData[43] ),
    .I1(\Inst_eFPGA_top.FrameData[44] ),
    .S(_0533_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1057_ (.I(_0537_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1058_ (.I(_0522_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1059_ (.I0(\Inst_eFPGA_top.FrameData[44] ),
    .I1(\Inst_eFPGA_top.FrameData[45] ),
    .S(_0538_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1060_ (.I(_0539_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1061_ (.I0(\Inst_eFPGA_top.FrameData[45] ),
    .I1(\Inst_eFPGA_top.FrameData[46] ),
    .S(_0538_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1062_ (.I(_0540_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1063_ (.I0(\Inst_eFPGA_top.FrameData[46] ),
    .I1(\Inst_eFPGA_top.FrameData[47] ),
    .S(_0538_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1064_ (.I(_0541_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1065_ (.I0(\Inst_eFPGA_top.FrameData[47] ),
    .I1(\Inst_eFPGA_top.FrameData[48] ),
    .S(_0538_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1066_ (.I(_0542_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1067_ (.I(_0521_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1068_ (.I(_0543_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1069_ (.I0(\Inst_eFPGA_top.FrameData[48] ),
    .I1(\Inst_eFPGA_top.FrameData[49] ),
    .S(_0544_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1070_ (.I(_0545_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1071_ (.I0(\Inst_eFPGA_top.FrameData[49] ),
    .I1(\Inst_eFPGA_top.FrameData[50] ),
    .S(_0544_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1072_ (.I(_0546_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1073_ (.I0(\Inst_eFPGA_top.FrameData[50] ),
    .I1(\Inst_eFPGA_top.FrameData[51] ),
    .S(_0544_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1074_ (.I(_0547_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1075_ (.I0(\Inst_eFPGA_top.FrameData[51] ),
    .I1(\Inst_eFPGA_top.FrameData[52] ),
    .S(_0544_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1076_ (.I(_0548_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1077_ (.I(_0543_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1078_ (.I0(\Inst_eFPGA_top.FrameData[52] ),
    .I1(\Inst_eFPGA_top.FrameData[53] ),
    .S(_0549_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1079_ (.I(_0550_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1080_ (.I0(\Inst_eFPGA_top.FrameData[53] ),
    .I1(\Inst_eFPGA_top.FrameData[54] ),
    .S(_0549_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1081_ (.I(_0551_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1082_ (.I0(\Inst_eFPGA_top.FrameData[54] ),
    .I1(\Inst_eFPGA_top.FrameData[55] ),
    .S(_0549_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1083_ (.I(_0552_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1084_ (.I0(\Inst_eFPGA_top.FrameData[55] ),
    .I1(\Inst_eFPGA_top.FrameData[56] ),
    .S(_0549_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1085_ (.I(_0553_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1086_ (.I(_0543_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1087_ (.I0(\Inst_eFPGA_top.FrameData[56] ),
    .I1(\Inst_eFPGA_top.FrameData[57] ),
    .S(_0554_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1088_ (.I(_0555_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1089_ (.I0(\Inst_eFPGA_top.FrameData[57] ),
    .I1(\Inst_eFPGA_top.FrameData[58] ),
    .S(_0554_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1090_ (.I(_0556_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1091_ (.I0(\Inst_eFPGA_top.FrameData[58] ),
    .I1(\Inst_eFPGA_top.FrameData[59] ),
    .S(_0554_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1092_ (.I(_0557_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1093_ (.I0(\Inst_eFPGA_top.FrameData[59] ),
    .I1(\Inst_eFPGA_top.FrameData[60] ),
    .S(_0554_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1094_ (.I(_0558_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1095_ (.I(_0543_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1096_ (.I0(\Inst_eFPGA_top.FrameData[60] ),
    .I1(\Inst_eFPGA_top.FrameData[61] ),
    .S(_0559_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1097_ (.I(_0560_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1098_ (.I0(\Inst_eFPGA_top.FrameData[61] ),
    .I1(\Inst_eFPGA_top.FrameData[62] ),
    .S(_0559_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1099_ (.I(_0561_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1100_ (.I0(\Inst_eFPGA_top.FrameData[62] ),
    .I1(\Inst_eFPGA_top.FrameData[63] ),
    .S(_0559_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1101_ (.I(_0562_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1102_ (.I0(\Inst_eFPGA_top.FrameData[63] ),
    .I1(\Inst_eFPGA_top.FrameData[64] ),
    .S(_0559_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1103_ (.I(_0563_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1104_ (.I(_0521_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1105_ (.I(_0564_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1106_ (.I0(\Inst_eFPGA_top.FrameData[64] ),
    .I1(\Inst_eFPGA_top.FrameData[65] ),
    .S(_0565_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1107_ (.I(_0566_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1108_ (.I0(\Inst_eFPGA_top.FrameData[65] ),
    .I1(\Inst_eFPGA_top.FrameData[66] ),
    .S(_0565_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1109_ (.I(_0567_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1110_ (.I0(\Inst_eFPGA_top.FrameData[66] ),
    .I1(\Inst_eFPGA_top.FrameData[67] ),
    .S(_0565_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1111_ (.I(_0568_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1112_ (.I0(\Inst_eFPGA_top.FrameData[67] ),
    .I1(\Inst_eFPGA_top.FrameData[68] ),
    .S(_0565_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1113_ (.I(_0569_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1114_ (.I(_0564_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1115_ (.I0(\Inst_eFPGA_top.FrameData[68] ),
    .I1(\Inst_eFPGA_top.FrameData[69] ),
    .S(_0570_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1116_ (.I(_0571_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1117_ (.I0(\Inst_eFPGA_top.FrameData[69] ),
    .I1(\Inst_eFPGA_top.FrameData[70] ),
    .S(_0570_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1118_ (.I(_0572_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1119_ (.I0(\Inst_eFPGA_top.FrameData[70] ),
    .I1(\Inst_eFPGA_top.FrameData[71] ),
    .S(_0570_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1120_ (.I(_0573_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1121_ (.I0(\Inst_eFPGA_top.FrameData[71] ),
    .I1(\Inst_eFPGA_top.FrameData[72] ),
    .S(_0570_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1122_ (.I(_0574_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1123_ (.I(_0564_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1124_ (.I0(\Inst_eFPGA_top.FrameData[72] ),
    .I1(\Inst_eFPGA_top.FrameData[73] ),
    .S(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1125_ (.I(_0576_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1126_ (.I0(\Inst_eFPGA_top.FrameData[73] ),
    .I1(\Inst_eFPGA_top.FrameData[74] ),
    .S(_0575_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1127_ (.I(_0577_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1128_ (.I0(\Inst_eFPGA_top.FrameData[74] ),
    .I1(\Inst_eFPGA_top.FrameData[75] ),
    .S(_0575_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1129_ (.I(_0578_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1130_ (.I0(\Inst_eFPGA_top.FrameData[75] ),
    .I1(\Inst_eFPGA_top.FrameData[76] ),
    .S(_0575_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1131_ (.I(_0579_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1132_ (.I(_0564_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1133_ (.I0(\Inst_eFPGA_top.FrameData[76] ),
    .I1(\Inst_eFPGA_top.FrameData[77] ),
    .S(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1134_ (.I(_0581_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1135_ (.I0(\Inst_eFPGA_top.FrameData[77] ),
    .I1(\Inst_eFPGA_top.FrameData[78] ),
    .S(_0580_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1136_ (.I(_0582_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1137_ (.I0(\Inst_eFPGA_top.FrameData[78] ),
    .I1(\Inst_eFPGA_top.FrameData[79] ),
    .S(_0580_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1138_ (.I(_0583_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1139_ (.I0(\Inst_eFPGA_top.FrameData[79] ),
    .I1(\Inst_eFPGA_top.FrameData[80] ),
    .S(_0580_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1140_ (.I(_0584_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1141_ (.I(_0521_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1142_ (.I(_0585_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1143_ (.I0(\Inst_eFPGA_top.FrameData[80] ),
    .I1(\Inst_eFPGA_top.FrameData[81] ),
    .S(_0586_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1144_ (.I(_0587_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1145_ (.I0(\Inst_eFPGA_top.FrameData[81] ),
    .I1(\Inst_eFPGA_top.FrameData[82] ),
    .S(_0586_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1146_ (.I(_0588_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1147_ (.I0(\Inst_eFPGA_top.FrameData[82] ),
    .I1(\Inst_eFPGA_top.FrameData[83] ),
    .S(_0586_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1148_ (.I(_0589_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1149_ (.I0(\Inst_eFPGA_top.FrameData[83] ),
    .I1(\Inst_eFPGA_top.FrameData[84] ),
    .S(_0586_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1150_ (.I(_0590_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1151_ (.I(_0585_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1152_ (.I0(\Inst_eFPGA_top.FrameData[84] ),
    .I1(\Inst_eFPGA_top.FrameData[85] ),
    .S(_0591_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1153_ (.I(_0592_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1154_ (.I0(\Inst_eFPGA_top.FrameData[85] ),
    .I1(\Inst_eFPGA_top.FrameData[86] ),
    .S(_0591_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1155_ (.I(_0593_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1156_ (.I0(\Inst_eFPGA_top.FrameData[86] ),
    .I1(\Inst_eFPGA_top.FrameData[87] ),
    .S(_0591_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1157_ (.I(_0594_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1158_ (.I0(\Inst_eFPGA_top.FrameData[87] ),
    .I1(\Inst_eFPGA_top.FrameData[88] ),
    .S(_0591_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1159_ (.I(_0595_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1160_ (.I(_0585_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1161_ (.I0(\Inst_eFPGA_top.FrameData[88] ),
    .I1(\Inst_eFPGA_top.FrameData[89] ),
    .S(_0596_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1162_ (.I(_0597_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1163_ (.I0(\Inst_eFPGA_top.FrameData[89] ),
    .I1(\Inst_eFPGA_top.FrameData[90] ),
    .S(_0596_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1164_ (.I(_0598_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1165_ (.I0(\Inst_eFPGA_top.FrameData[90] ),
    .I1(\Inst_eFPGA_top.FrameData[91] ),
    .S(_0596_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1166_ (.I(_0599_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1167_ (.I0(\Inst_eFPGA_top.FrameData[91] ),
    .I1(\Inst_eFPGA_top.FrameData[92] ),
    .S(_0596_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1168_ (.I(_0600_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1169_ (.I(_0585_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1170_ (.I0(\Inst_eFPGA_top.FrameData[92] ),
    .I1(\Inst_eFPGA_top.FrameData[93] ),
    .S(_0601_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1171_ (.I(_0602_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1172_ (.I0(\Inst_eFPGA_top.FrameData[93] ),
    .I1(\Inst_eFPGA_top.FrameData[94] ),
    .S(_0601_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1173_ (.I(_0603_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1174_ (.I0(\Inst_eFPGA_top.FrameData[94] ),
    .I1(\Inst_eFPGA_top.FrameData[95] ),
    .S(_0601_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1175_ (.I(_0604_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1176_ (.I0(\Inst_eFPGA_top.FrameData[95] ),
    .I1(\Inst_eFPGA_top.FrameData[96] ),
    .S(_0601_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1177_ (.I(_0605_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1178_ (.I(net18),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1179_ (.I(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1180_ (.I0(\Inst_eFPGA_top.FrameData[96] ),
    .I1(\Inst_eFPGA_top.FrameData[97] ),
    .S(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1181_ (.I(_0608_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1182_ (.I0(\Inst_eFPGA_top.FrameData[97] ),
    .I1(\Inst_eFPGA_top.FrameData[98] ),
    .S(_0607_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1183_ (.I(_0609_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1184_ (.I0(\Inst_eFPGA_top.FrameData[98] ),
    .I1(\Inst_eFPGA_top.FrameData[99] ),
    .S(_0607_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1185_ (.I(_0610_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1186_ (.I0(\Inst_eFPGA_top.FrameData[99] ),
    .I1(\Inst_eFPGA_top.FrameData[100] ),
    .S(_0607_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1187_ (.I(_0611_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1188_ (.I(_0606_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1189_ (.I0(\Inst_eFPGA_top.FrameData[100] ),
    .I1(\Inst_eFPGA_top.FrameData[101] ),
    .S(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1190_ (.I(_0613_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1191_ (.I0(\Inst_eFPGA_top.FrameData[101] ),
    .I1(\Inst_eFPGA_top.FrameData[102] ),
    .S(_0612_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1192_ (.I(_0614_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1193_ (.I0(\Inst_eFPGA_top.FrameData[102] ),
    .I1(\Inst_eFPGA_top.FrameData[103] ),
    .S(_0612_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1194_ (.I(_0615_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1195_ (.I0(\Inst_eFPGA_top.FrameData[103] ),
    .I1(\Inst_eFPGA_top.FrameData[104] ),
    .S(_0612_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1196_ (.I(_0616_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1197_ (.I(_0606_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1198_ (.I0(\Inst_eFPGA_top.FrameData[104] ),
    .I1(\Inst_eFPGA_top.FrameData[105] ),
    .S(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1199_ (.I(_0618_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1200_ (.I0(\Inst_eFPGA_top.FrameData[105] ),
    .I1(\Inst_eFPGA_top.FrameData[106] ),
    .S(_0617_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1201_ (.I(_0619_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1202_ (.I0(\Inst_eFPGA_top.FrameData[106] ),
    .I1(\Inst_eFPGA_top.FrameData[107] ),
    .S(_0617_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1203_ (.I(_0620_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1204_ (.I0(\Inst_eFPGA_top.FrameData[107] ),
    .I1(\Inst_eFPGA_top.FrameData[108] ),
    .S(_0617_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1205_ (.I(_0621_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1206_ (.I(_0606_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1207_ (.I0(\Inst_eFPGA_top.FrameData[108] ),
    .I1(\Inst_eFPGA_top.FrameData[109] ),
    .S(_0622_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1208_ (.I(_0623_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1209_ (.I0(\Inst_eFPGA_top.FrameData[109] ),
    .I1(\Inst_eFPGA_top.FrameData[110] ),
    .S(_0622_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1210_ (.I(_0624_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1211_ (.I0(\Inst_eFPGA_top.FrameData[110] ),
    .I1(\Inst_eFPGA_top.FrameData[111] ),
    .S(_0622_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1212_ (.I(_0625_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1213_ (.I0(\Inst_eFPGA_top.FrameData[111] ),
    .I1(\Inst_eFPGA_top.FrameData[112] ),
    .S(_0622_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1214_ (.I(_0294_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1215_ (.I(net18),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1216_ (.I(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1217_ (.I0(\Inst_eFPGA_top.FrameData[112] ),
    .I1(\Inst_eFPGA_top.FrameData[113] ),
    .S(_0296_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1218_ (.I(_0297_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1219_ (.I0(\Inst_eFPGA_top.FrameData[113] ),
    .I1(\Inst_eFPGA_top.FrameData[114] ),
    .S(_0296_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1220_ (.I(_0298_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1221_ (.I0(\Inst_eFPGA_top.FrameData[114] ),
    .I1(\Inst_eFPGA_top.FrameData[115] ),
    .S(_0296_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1222_ (.I(_0299_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1223_ (.I0(\Inst_eFPGA_top.FrameData[115] ),
    .I1(\Inst_eFPGA_top.FrameData[116] ),
    .S(_0296_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1224_ (.I(_0300_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1225_ (.I(_0295_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1226_ (.I0(\Inst_eFPGA_top.FrameData[116] ),
    .I1(\Inst_eFPGA_top.FrameData[117] ),
    .S(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1227_ (.I(_0302_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1228_ (.I0(\Inst_eFPGA_top.FrameData[117] ),
    .I1(\Inst_eFPGA_top.FrameData[118] ),
    .S(_0301_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1229_ (.I(_0303_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1230_ (.I0(\Inst_eFPGA_top.FrameData[118] ),
    .I1(\Inst_eFPGA_top.FrameData[119] ),
    .S(_0301_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1231_ (.I(_0304_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1232_ (.I0(\Inst_eFPGA_top.FrameData[119] ),
    .I1(\Inst_eFPGA_top.FrameData[120] ),
    .S(_0301_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1233_ (.I(_0305_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1234_ (.I(_0295_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1235_ (.I0(\Inst_eFPGA_top.FrameData[120] ),
    .I1(\Inst_eFPGA_top.FrameData[121] ),
    .S(_0306_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1236_ (.I(_0307_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1237_ (.I0(\Inst_eFPGA_top.FrameData[121] ),
    .I1(\Inst_eFPGA_top.FrameData[122] ),
    .S(_0306_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1238_ (.I(_0308_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1239_ (.I0(\Inst_eFPGA_top.FrameData[122] ),
    .I1(\Inst_eFPGA_top.FrameData[123] ),
    .S(_0306_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1240_ (.I(_0309_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1241_ (.I0(\Inst_eFPGA_top.FrameData[123] ),
    .I1(\Inst_eFPGA_top.FrameData[124] ),
    .S(_0306_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1242_ (.I(_0310_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _1243_ (.I(_0295_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1244_ (.I0(\Inst_eFPGA_top.FrameData[124] ),
    .I1(\Inst_eFPGA_top.FrameData[125] ),
    .S(_0311_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1245_ (.I(_0312_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1246_ (.I0(\Inst_eFPGA_top.FrameData[125] ),
    .I1(\Inst_eFPGA_top.FrameData[126] ),
    .S(_0311_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1247_ (.I(_0313_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1248_ (.I0(\Inst_eFPGA_top.FrameData[126] ),
    .I1(\Inst_eFPGA_top.FrameData[127] ),
    .S(_0311_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1249_ (.I(_0314_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1250_ (.I0(\Inst_eFPGA_top.FrameData[127] ),
    .I1(net19),
    .S(_0311_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1251_ (.I(_0315_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1252_ (.D(_0188_),
    .CLK(clknet_4_5_0_io_in[5]),
    .Q(\fstb_ctr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1253_ (.D(_0189_),
    .CLK(clknet_4_6_0_io_in[5]),
    .Q(\fstb_ctr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1254_ (.D(_0190_),
    .CLK(clknet_4_5_0_io_in[5]),
    .Q(\fstb_ctr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1255_ (.D(_0191_),
    .CLK(clknet_4_7_0_io_in[5]),
    .Q(\fstb_ctr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1256_ (.D(_0192_),
    .CLK(clknet_4_7_0_io_in[5]),
    .Q(\fstb_ctr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1257_ (.D(_0193_),
    .CLK(clknet_4_4_0_io_in[5]),
    .Q(\fstb_ctr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1258_ (.D(_0194_),
    .CLK(clknet_4_4_0_io_in[5]),
    .Q(\fstb_ctr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1259_ (.D(_0195_),
    .CLK(clknet_4_5_0_io_in[5]),
    .Q(\fstb_ctr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1260_ (.D(_0196_),
    .CLK(clknet_4_6_0_io_in[5]),
    .Q(\fstb_ctr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1261_ (.D(_0197_),
    .CLK(clknet_4_5_0_io_in[5]),
    .Q(\fstb_ctr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1262_ (.D(_0198_),
    .CLK(clknet_4_7_0_io_in[5]),
    .Q(\fstb_ctr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1263_ (.D(_0199_),
    .CLK(clknet_4_6_0_io_in[5]),
    .Q(\fstb_ctr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1264_ (.D(_0200_),
    .CLK(clknet_4_7_0_io_in[5]),
    .Q(\fstb_ctr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1265_ (.D(_0201_),
    .CLK(clknet_4_6_0_io_in[5]),
    .Q(\fstb_ctr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1266_ (.D(_0202_),
    .CLK(clknet_4_7_0_io_in[5]),
    .Q(\fstb_ctr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1267_ (.D(_0203_),
    .CLK(clknet_4_4_0_io_in[5]),
    .Q(\fstb_ctr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1268_ (.D(_0204_),
    .CLK(clknet_4_10_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1269_ (.D(_0205_),
    .CLK(clknet_4_10_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1270_ (.D(_0206_),
    .CLK(clknet_4_14_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1271_ (.D(_0207_),
    .CLK(clknet_4_14_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1272_ (.D(_0208_),
    .CLK(clknet_4_10_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1273_ (.D(_0209_),
    .CLK(clknet_4_11_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1274_ (.D(_0210_),
    .CLK(clknet_4_14_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1275_ (.D(_0211_),
    .CLK(clknet_4_10_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1276_ (.D(_0212_),
    .CLK(clknet_4_14_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1277_ (.D(_0213_),
    .CLK(clknet_4_8_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1278_ (.D(_0214_),
    .CLK(clknet_4_8_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1279_ (.D(_0215_),
    .CLK(clknet_4_8_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1280_ (.D(_0216_),
    .CLK(clknet_4_8_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1281_ (.D(_0217_),
    .CLK(clknet_4_10_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1282_ (.D(_0218_),
    .CLK(clknet_4_8_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1283_ (.D(_0219_),
    .CLK(clknet_4_10_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1284_ (.D(_0220_),
    .CLK(clknet_4_10_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1285_ (.D(_0221_),
    .CLK(clknet_4_14_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1286_ (.D(_0222_),
    .CLK(clknet_4_8_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1287_ (.D(_0223_),
    .CLK(clknet_4_11_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1288_ (.D(_0224_),
    .CLK(clknet_4_14_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1289_ (.D(_0225_),
    .CLK(clknet_4_11_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1290_ (.D(_0226_),
    .CLK(clknet_4_11_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1291_ (.D(_0227_),
    .CLK(clknet_4_11_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1292_ (.D(_0228_),
    .CLK(clknet_4_11_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1293_ (.D(_0229_),
    .CLK(clknet_4_11_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1294_ (.D(_0230_),
    .CLK(clknet_4_11_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1295_ (.D(_0231_),
    .CLK(clknet_4_14_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1296_ (.D(_0232_),
    .CLK(clknet_4_14_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1297_ (.D(_0233_),
    .CLK(clknet_4_14_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1298_ (.D(_0234_),
    .CLK(clknet_4_11_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1299_ (.D(_0235_),
    .CLK(clknet_4_8_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1300_ (.D(_0236_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[64] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1301_ (.D(_0237_),
    .CLK(clknet_4_13_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[65] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1302_ (.D(_0238_),
    .CLK(clknet_4_13_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[66] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1303_ (.D(_0239_),
    .CLK(clknet_4_13_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[67] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1304_ (.D(_0240_),
    .CLK(clknet_4_13_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[68] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1305_ (.D(_0241_),
    .CLK(clknet_4_13_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[69] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1306_ (.D(_0242_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[70] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1307_ (.D(_0243_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[71] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1308_ (.D(_0244_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[72] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1309_ (.D(_0245_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[73] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1310_ (.D(_0246_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[74] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1311_ (.D(_0247_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[75] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1312_ (.D(_0248_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[76] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1313_ (.D(_0249_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[77] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1314_ (.D(_0250_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[78] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1315_ (.D(_0251_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[79] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1316_ (.D(_0252_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[80] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1317_ (.D(_0253_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[81] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1318_ (.D(_0254_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[82] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1319_ (.D(_0255_),
    .CLK(clknet_4_15_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[83] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1320_ (.D(_0256_),
    .CLK(clknet_4_15_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[84] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1321_ (.D(_0257_),
    .CLK(clknet_4_15_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[85] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1322_ (.D(_0258_),
    .CLK(clknet_4_15_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[86] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1323_ (.D(_0259_),
    .CLK(clknet_4_15_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[87] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1324_ (.D(_0260_),
    .CLK(clknet_4_9_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[88] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1325_ (.D(_0261_),
    .CLK(clknet_4_9_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[89] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1326_ (.D(_0262_),
    .CLK(clknet_4_9_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[90] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1327_ (.D(_0263_),
    .CLK(clknet_4_9_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[91] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1328_ (.D(_0264_),
    .CLK(clknet_4_15_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[92] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1329_ (.D(_0265_),
    .CLK(clknet_4_9_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[93] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1330_ (.D(_0266_),
    .CLK(clknet_4_15_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[94] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1331_ (.D(_0267_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[95] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1332_ (.D(_0268_),
    .CLK(clknet_4_3_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[96] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1333_ (.D(_0269_),
    .CLK(clknet_4_0_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[97] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1334_ (.D(_0270_),
    .CLK(clknet_4_0_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[98] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1335_ (.D(_0271_),
    .CLK(clknet_4_0_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[99] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1336_ (.D(_0272_),
    .CLK(clknet_4_0_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[100] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1337_ (.D(_0273_),
    .CLK(clknet_4_0_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[101] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1338_ (.D(_0274_),
    .CLK(clknet_4_1_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[102] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1339_ (.D(_0275_),
    .CLK(clknet_4_1_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[103] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1340_ (.D(_0276_),
    .CLK(clknet_4_1_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[104] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1341_ (.D(_0277_),
    .CLK(clknet_4_1_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[105] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1342_ (.D(_0278_),
    .CLK(clknet_4_1_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[106] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1343_ (.D(_0279_),
    .CLK(clknet_4_1_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[107] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1344_ (.D(_0280_),
    .CLK(clknet_4_3_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[108] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1345_ (.D(_0281_),
    .CLK(clknet_4_1_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[109] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1346_ (.D(_0282_),
    .CLK(clknet_4_3_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[110] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1347_ (.D(_0283_),
    .CLK(clknet_4_3_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[111] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1348_ (.D(_0284_),
    .CLK(clknet_4_3_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[112] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1349_ (.D(_0285_),
    .CLK(clknet_4_3_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[113] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1350_ (.D(_0286_),
    .CLK(clknet_4_2_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[114] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1351_ (.D(_0287_),
    .CLK(clknet_4_2_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[115] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1352_ (.D(_0288_),
    .CLK(clknet_4_2_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[116] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1353_ (.D(_0289_),
    .CLK(clknet_4_2_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[117] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1354_ (.D(_0290_),
    .CLK(clknet_4_2_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[118] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1355_ (.D(_0291_),
    .CLK(clknet_4_2_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[119] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1356_ (.D(_0292_),
    .CLK(clknet_4_2_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[120] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1357_ (.D(_0293_),
    .CLK(clknet_4_2_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[121] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1358_ (.D(_0182_),
    .CLK(clknet_4_2_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[122] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1359_ (.D(_0183_),
    .CLK(clknet_4_13_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[123] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1360_ (.D(_0184_),
    .CLK(clknet_4_13_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[124] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1361_ (.D(_0185_),
    .CLK(clknet_4_13_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[125] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1362_ (.D(_0186_),
    .CLK(clknet_4_13_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[126] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1363_ (.D(_0187_),
    .CLK(clknet_4_12_0_io_in[5]),
    .Q(\Inst_eFPGA_top.FrameData[127] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_186 (.Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_187 (.Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_188 (.Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_189 (.Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_190 (.Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_191 (.Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_192 (.Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_193 (.Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_194 (.Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_195 (.Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_0_io_in[5]  (.I(io_in[5]),
    .Z(clknet_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_example_185 (.Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1509_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_T_top ),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1510_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_T_top ),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1511_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_T_top ),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1512_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_T_top ),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1513_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_T_top ),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1514_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_T_top ),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1515_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_T_top ),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1516_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_T_top ),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1517_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_T_top ),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1518_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_T_top ),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1519_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_T_top ),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1520_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_T_top ),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1521_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_I_top ),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1522_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_I_top ),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1523_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_I_top ),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1524_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_I_top ),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1525_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_I_top ),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1526_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_I_top ),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1527_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_I_top ),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1528_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_I_top ),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1529_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_I_top ),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1530_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_I_top ),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1531_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_I_top ),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1532_ (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_I_top ),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[0].rs_and  (.A1(_0040_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[100].rs_and  (.A1(_0013_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[100] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[101].rs_and  (.A1(_0014_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[101] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[102].rs_and  (.A1(_0015_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[102] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[103].rs_and  (.A1(_0016_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[103] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[104].rs_and  (.A1(_0017_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[104] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[105].rs_and  (.A1(_0018_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[105] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[106].rs_and  (.A1(_0019_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[106] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[107].rs_and  (.A1(_0020_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[107] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[108].rs_and  (.A1(_0021_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[108] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[109].rs_and  (.A1(_0022_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[109] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[10].rs_and  (.A1(_0103_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[10] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[110].rs_and  (.A1(_0023_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[110] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[111].rs_and  (.A1(_0024_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[111] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[112].rs_and  (.A1(_0025_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[112] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[113].rs_and  (.A1(_0026_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[113] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[114].rs_and  (.A1(_0027_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[114] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[115].rs_and  (.A1(_0028_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[115] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[116].rs_and  (.A1(_0029_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[116] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[117].rs_and  (.A1(_0030_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[117] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[118].rs_and  (.A1(_0031_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[118] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[119].rs_and  (.A1(_0032_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[119] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[11].rs_and  (.A1(_0104_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[11] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[120].rs_and  (.A1(_0033_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[120] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[121].rs_and  (.A1(_0034_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[121] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[122].rs_and  (.A1(_0035_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[122] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[123].rs_and  (.A1(_0036_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[123] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[124].rs_and  (.A1(_0037_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[124] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[125].rs_and  (.A1(_0038_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[125] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[126].rs_and  (.A1(_0039_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[126] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[127].rs_and  (.A1(_0041_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[127] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[128].rs_and  (.A1(_0042_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[128] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[129].rs_and  (.A1(_0043_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[129] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[12].rs_and  (.A1(_0105_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[12] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[130].rs_and  (.A1(_0044_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[130] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[131].rs_and  (.A1(_0045_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[131] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[132].rs_and  (.A1(_0046_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[132] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[133].rs_and  (.A1(_0047_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[133] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[134].rs_and  (.A1(_0048_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[134] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[135].rs_and  (.A1(_0049_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[135] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[136].rs_and  (.A1(_0050_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[136] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[137].rs_and  (.A1(_0052_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[137] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[138].rs_and  (.A1(_0053_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[138] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[139].rs_and  (.A1(_0054_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[139] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[13].rs_and  (.A1(_0106_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[13] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[140].rs_and  (.A1(_0055_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[140] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[141].rs_and  (.A1(_0056_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[141] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[142].rs_and  (.A1(_0057_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[142] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[143].rs_and  (.A1(_0058_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[143] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[144].rs_and  (.A1(_0059_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[144] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[145].rs_and  (.A1(_0060_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[145] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[146].rs_and  (.A1(_0061_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[146] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[147].rs_and  (.A1(_0063_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[147] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[148].rs_and  (.A1(_0064_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[148] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[149].rs_and  (.A1(_0065_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[149] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[14].rs_and  (.A1(_0107_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[14] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[150].rs_and  (.A1(_0066_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[150] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[151].rs_and  (.A1(_0067_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[151] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[152].rs_and  (.A1(_0068_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[152] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[153].rs_and  (.A1(_0069_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[153] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[154].rs_and  (.A1(_0070_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[154] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[155].rs_and  (.A1(_0071_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[155] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[156].rs_and  (.A1(_0072_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[156] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[157].rs_and  (.A1(_0074_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[157] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[158].rs_and  (.A1(_0075_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[158] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[159].rs_and  (.A1(_0076_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[159] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[15].rs_and  (.A1(_0108_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[15] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[160].rs_and  (.A1(_0077_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[160] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[161].rs_and  (.A1(_0078_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[161] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[162].rs_and  (.A1(_0079_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[162] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[163].rs_and  (.A1(_0080_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[163] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[164].rs_and  (.A1(_0081_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[164] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[165].rs_and  (.A1(_0082_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[165] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[166].rs_and  (.A1(_0083_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[166] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[167].rs_and  (.A1(_0085_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[167] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[168].rs_and  (.A1(_0086_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[168] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[169].rs_and  (.A1(_0087_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[169] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[16].rs_and  (.A1(_0109_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[16] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[170].rs_and  (.A1(_0088_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[170] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[171].rs_and  (.A1(_0089_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[171] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[172].rs_and  (.A1(_0090_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[172] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[173].rs_and  (.A1(_0091_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[173] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[174].rs_and  (.A1(_0092_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[174] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[175].rs_and  (.A1(_0093_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[175] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[176].rs_and  (.A1(_0094_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[176] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[177].rs_and  (.A1(_0096_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[177] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[178].rs_and  (.A1(_0097_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[178] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[179].rs_and  (.A1(_0098_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[179] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[17].rs_and  (.A1(_0110_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[17] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[18].rs_and  (.A1(_0111_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[18] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[19].rs_and  (.A1(_0112_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[19] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[1].rs_and  (.A1(_0051_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[1] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[20].rs_and  (.A1(_0113_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[20] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[21].rs_and  (.A1(_0114_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[21] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[22].rs_and  (.A1(_0115_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[22] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[23].rs_and  (.A1(_0116_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[23] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[24].rs_and  (.A1(_0117_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[24] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[25].rs_and  (.A1(_0118_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[25] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[26].rs_and  (.A1(_0119_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[26] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[27].rs_and  (.A1(_0120_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[27] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[28].rs_and  (.A1(_0121_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[28] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[29].rs_and  (.A1(_0122_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[29] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[2].rs_and  (.A1(_0062_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[2] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[30].rs_and  (.A1(_0123_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[30] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[31].rs_and  (.A1(_0124_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[31] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[32].rs_and  (.A1(_0125_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[32] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[33].rs_and  (.A1(_0126_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[33] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[34].rs_and  (.A1(_0127_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[34] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[35].rs_and  (.A1(_0128_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[35] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[36].rs_and  (.A1(_0129_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[36] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[37].rs_and  (.A1(_0130_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[37] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[38].rs_and  (.A1(_0131_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[38] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[39].rs_and  (.A1(_0132_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[39] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[3].rs_and  (.A1(_0073_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[3] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[40].rs_and  (.A1(_0133_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[40] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[41].rs_and  (.A1(_0134_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[41] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[42].rs_and  (.A1(_0135_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[42] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[43].rs_and  (.A1(_0136_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[43] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[44].rs_and  (.A1(_0137_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[44] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[45].rs_and  (.A1(_0138_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[45] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[46].rs_and  (.A1(_0139_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[46] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[47].rs_and  (.A1(_0140_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[47] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[48].rs_and  (.A1(_0141_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[48] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[49].rs_and  (.A1(_0142_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[49] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[4].rs_and  (.A1(_0084_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[4] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[50].rs_and  (.A1(_0143_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[50] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[51].rs_and  (.A1(_0144_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[51] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[52].rs_and  (.A1(_0145_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[52] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[53].rs_and  (.A1(_0146_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[53] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[54].rs_and  (.A1(_0147_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[54] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[55].rs_and  (.A1(_0148_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[55] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[56].rs_and  (.A1(_0149_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[56] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[57].rs_and  (.A1(_0150_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[57] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[58].rs_and  (.A1(_0151_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[58] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[59].rs_and  (.A1(_0152_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[59] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[5].rs_and  (.A1(_0095_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[5] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[60].rs_and  (.A1(_0153_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[60] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[61].rs_and  (.A1(_0154_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[61] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[62].rs_and  (.A1(_0155_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[62] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[63].rs_and  (.A1(_0156_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[63] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[64].rs_and  (.A1(_0157_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[64] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[65].rs_and  (.A1(_0158_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[65] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[66].rs_and  (.A1(_0159_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[66] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[67].rs_and  (.A1(_0160_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[67] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[68].rs_and  (.A1(_0161_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[68] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[69].rs_and  (.A1(_0162_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[69] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[6].rs_and  (.A1(_0099_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[6] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[70].rs_and  (.A1(_0163_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[70] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[71].rs_and  (.A1(_0164_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[71] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[72].rs_and  (.A1(_0165_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[72] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[73].rs_and  (.A1(_0166_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[73] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[74].rs_and  (.A1(_0167_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[74] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[75].rs_and  (.A1(_0168_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[75] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[76].rs_and  (.A1(_0169_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[76] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[77].rs_and  (.A1(_0170_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[77] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[78].rs_and  (.A1(_0171_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[78] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[79].rs_and  (.A1(_0172_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[79] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[7].rs_and  (.A1(_0100_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[7] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[80].rs_and  (.A1(_0173_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[80] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[81].rs_and  (.A1(_0174_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[81] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[82].rs_and  (.A1(_0175_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[82] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[83].rs_and  (.A1(_0176_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[83] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[84].rs_and  (.A1(_0177_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[84] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[85].rs_and  (.A1(_0178_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[85] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[86].rs_and  (.A1(_0179_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[86] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[87].rs_and  (.A1(_0000_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[87] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[88].rs_and  (.A1(_0001_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[88] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[89].rs_and  (.A1(_0002_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[89] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[8].rs_and  (.A1(_0101_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[8] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[90].rs_and  (.A1(_0003_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[90] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[91].rs_and  (.A1(_0004_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[91] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[92].rs_and  (.A1(_0005_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[92] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[93].rs_and  (.A1(_0006_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[93] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[94].rs_and  (.A1(_0007_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[94] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[95].rs_and  (.A1(_0008_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[95] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[96].rs_and  (.A1(_0009_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[96] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[97].rs_and  (.A1(_0010_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[97] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[98].rs_and  (.A1(_0011_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[98] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[99].rs_and  (.A1(_0012_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[99] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \frame_ands[9].rs_and  (.A1(_0102_),
    .A2(net1),
    .Z(\Inst_eFPGA_top.FrameSelect[9] ));
 gf180mcu_fpga_bitmux sram_test0_i (.BLP(net4),
    .BLN(_0180_),
    .WL(net3),
    .I(net22),
    .O(net48));
 gf180mcu_fpga_bitmux sram_test1_i (.BLP(net5),
    .BLN(_0181_),
    .WL(net3),
    .I(net23),
    .O(net49));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[16]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[17]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[18]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(io_in[26]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[27]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input8 (.I(io_in[28]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(io_in[29]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(io_in[30]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(io_in[31]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input12 (.I(io_in[32]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input13 (.I(io_in[33]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(io_in[34]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(io_in[35]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input16 (.I(io_in[36]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input17 (.I(io_in[37]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(io_in[6]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(io_in[7]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input20 (.I(io_in[8]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input21 (.I(io_in[9]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(la_data_in[0]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(la_data_in[1]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output24 (.I(net24),
    .Z(io_oeb[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output25 (.I(net25),
    .Z(io_oeb[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output26 (.I(net26),
    .Z(io_oeb[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output27 (.I(net27),
    .Z(io_oeb[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output28 (.I(net28),
    .Z(io_oeb[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output29 (.I(net29),
    .Z(io_oeb[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output30 (.I(net30),
    .Z(io_oeb[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output31 (.I(net31),
    .Z(io_oeb[33]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output32 (.I(net32),
    .Z(io_oeb[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output33 (.I(net33),
    .Z(io_oeb[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output34 (.I(net34),
    .Z(io_oeb[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output35 (.I(net35),
    .Z(io_oeb[37]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output36 (.I(net36),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output37 (.I(net37),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output38 (.I(net38),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output39 (.I(net39),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output40 (.I(net40),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output41 (.I(net41),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output42 (.I(net42),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output43 (.I(net43),
    .Z(io_out[33]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output44 (.I(net44),
    .Z(io_out[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output45 (.I(net45),
    .Z(io_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output46 (.I(net46),
    .Z(io_out[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output47 (.I(net47),
    .Z(io_out[37]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output48 (.I(net48),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output49 (.I(net49),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout50 (.I(net2),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_example_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_2_0_0_io_in[5]  (.I(clknet_0_io_in[5]),
    .Z(clknet_2_0_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_2_1_0_io_in[5]  (.I(clknet_0_io_in[5]),
    .Z(clknet_2_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_2_2_0_io_in[5]  (.I(clknet_0_io_in[5]),
    .Z(clknet_2_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_2_3_0_io_in[5]  (.I(clknet_0_io_in[5]),
    .Z(clknet_2_3_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_0_0_io_in[5]  (.I(clknet_2_0_0_io_in[5]),
    .Z(clknet_3_0_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_0_1_io_in[5]  (.I(clknet_3_0_0_io_in[5]),
    .Z(clknet_3_0_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_1_0_io_in[5]  (.I(clknet_2_0_0_io_in[5]),
    .Z(clknet_3_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_1_1_io_in[5]  (.I(clknet_3_1_0_io_in[5]),
    .Z(clknet_3_1_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_2_0_io_in[5]  (.I(clknet_2_1_0_io_in[5]),
    .Z(clknet_3_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_2_1_io_in[5]  (.I(clknet_3_2_0_io_in[5]),
    .Z(clknet_3_2_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_3_0_io_in[5]  (.I(clknet_2_1_0_io_in[5]),
    .Z(clknet_3_3_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_3_1_io_in[5]  (.I(clknet_3_3_0_io_in[5]),
    .Z(clknet_3_3_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_4_0_io_in[5]  (.I(clknet_2_2_0_io_in[5]),
    .Z(clknet_3_4_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_4_1_io_in[5]  (.I(clknet_3_4_0_io_in[5]),
    .Z(clknet_3_4_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_5_0_io_in[5]  (.I(clknet_2_2_0_io_in[5]),
    .Z(clknet_3_5_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_5_1_io_in[5]  (.I(clknet_3_5_0_io_in[5]),
    .Z(clknet_3_5_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_6_0_io_in[5]  (.I(clknet_2_3_0_io_in[5]),
    .Z(clknet_3_6_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_6_1_io_in[5]  (.I(clknet_3_6_0_io_in[5]),
    .Z(clknet_3_6_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_7_0_io_in[5]  (.I(clknet_2_3_0_io_in[5]),
    .Z(clknet_3_7_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_3_7_1_io_in[5]  (.I(clknet_3_7_0_io_in[5]),
    .Z(clknet_3_7_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_0_0_io_in[5]  (.I(clknet_3_0_1_io_in[5]),
    .Z(clknet_4_0_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_1_0_io_in[5]  (.I(clknet_3_0_1_io_in[5]),
    .Z(clknet_4_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_2_0_io_in[5]  (.I(clknet_3_1_1_io_in[5]),
    .Z(clknet_4_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_3_0_io_in[5]  (.I(clknet_3_1_1_io_in[5]),
    .Z(clknet_4_3_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_4_0_io_in[5]  (.I(clknet_3_2_1_io_in[5]),
    .Z(clknet_4_4_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_5_0_io_in[5]  (.I(clknet_3_2_1_io_in[5]),
    .Z(clknet_4_5_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_6_0_io_in[5]  (.I(clknet_3_3_1_io_in[5]),
    .Z(clknet_4_6_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_7_0_io_in[5]  (.I(clknet_3_3_1_io_in[5]),
    .Z(clknet_4_7_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_8_0_io_in[5]  (.I(clknet_3_4_1_io_in[5]),
    .Z(clknet_4_8_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_9_0_io_in[5]  (.I(clknet_3_4_1_io_in[5]),
    .Z(clknet_4_9_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_10_0_io_in[5]  (.I(clknet_3_5_1_io_in[5]),
    .Z(clknet_4_10_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_11_0_io_in[5]  (.I(clknet_3_5_1_io_in[5]),
    .Z(clknet_4_11_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_12_0_io_in[5]  (.I(clknet_3_6_1_io_in[5]),
    .Z(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_13_0_io_in[5]  (.I(clknet_3_6_1_io_in[5]),
    .Z(clknet_4_13_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_14_0_io_in[5]  (.I(clknet_3_7_1_io_in[5]),
    .Z(clknet_4_14_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \clkbuf_4_15_0_io_in[5]  (.I(clknet_3_7_1_io_in[5]),
    .Z(clknet_4_15_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_opt_1_0_io_in[5]  (.I(clknet_4_7_0_io_in[5]),
    .Z(clknet_opt_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_opt_1_1_io_in[5]  (.I(clknet_opt_1_0_io_in[5]),
    .Z(clknet_opt_1_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_opt_1_2_io_in[5]  (.I(clknet_opt_1_1_io_in[5]),
    .Z(clknet_opt_1_2_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1189__I0 (.I(\Inst_eFPGA_top.FrameData[100] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1186__I1 (.I(\Inst_eFPGA_top.FrameData[100] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[4]  (.I(\Inst_eFPGA_top.FrameData[100] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1191__I0 (.I(\Inst_eFPGA_top.FrameData[101] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1189__I1 (.I(\Inst_eFPGA_top.FrameData[101] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[5]  (.I(\Inst_eFPGA_top.FrameData[101] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1193__I0 (.I(\Inst_eFPGA_top.FrameData[102] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1191__I1 (.I(\Inst_eFPGA_top.FrameData[102] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[6]  (.I(\Inst_eFPGA_top.FrameData[102] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1207__I0 (.I(\Inst_eFPGA_top.FrameData[108] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1204__I1 (.I(\Inst_eFPGA_top.FrameData[108] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[12]  (.I(\Inst_eFPGA_top.FrameData[108] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1211__I0 (.I(\Inst_eFPGA_top.FrameData[110] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1209__I1 (.I(\Inst_eFPGA_top.FrameData[110] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[14]  (.I(\Inst_eFPGA_top.FrameData[110] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1217__I0 (.I(\Inst_eFPGA_top.FrameData[112] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1213__I1 (.I(\Inst_eFPGA_top.FrameData[112] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[16]  (.I(\Inst_eFPGA_top.FrameData[112] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1221__I0 (.I(\Inst_eFPGA_top.FrameData[114] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1219__I1 (.I(\Inst_eFPGA_top.FrameData[114] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[18]  (.I(\Inst_eFPGA_top.FrameData[114] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1223__I0 (.I(\Inst_eFPGA_top.FrameData[115] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1221__I1 (.I(\Inst_eFPGA_top.FrameData[115] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[19]  (.I(\Inst_eFPGA_top.FrameData[115] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1226__I0 (.I(\Inst_eFPGA_top.FrameData[116] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1223__I1 (.I(\Inst_eFPGA_top.FrameData[116] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[20]  (.I(\Inst_eFPGA_top.FrameData[116] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1228__I0 (.I(\Inst_eFPGA_top.FrameData[117] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1226__I1 (.I(\Inst_eFPGA_top.FrameData[117] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[21]  (.I(\Inst_eFPGA_top.FrameData[117] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1230__I0 (.I(\Inst_eFPGA_top.FrameData[118] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1228__I1 (.I(\Inst_eFPGA_top.FrameData[118] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[22]  (.I(\Inst_eFPGA_top.FrameData[118] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1232__I0 (.I(\Inst_eFPGA_top.FrameData[119] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1230__I1 (.I(\Inst_eFPGA_top.FrameData[119] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[23]  (.I(\Inst_eFPGA_top.FrameData[119] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1235__I0 (.I(\Inst_eFPGA_top.FrameData[120] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1232__I1 (.I(\Inst_eFPGA_top.FrameData[120] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[24]  (.I(\Inst_eFPGA_top.FrameData[120] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1237__I0 (.I(\Inst_eFPGA_top.FrameData[121] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1235__I1 (.I(\Inst_eFPGA_top.FrameData[121] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[25]  (.I(\Inst_eFPGA_top.FrameData[121] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1239__I0 (.I(\Inst_eFPGA_top.FrameData[122] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1237__I1 (.I(\Inst_eFPGA_top.FrameData[122] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[26]  (.I(\Inst_eFPGA_top.FrameData[122] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1241__I0 (.I(\Inst_eFPGA_top.FrameData[123] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1239__I1 (.I(\Inst_eFPGA_top.FrameData[123] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[27]  (.I(\Inst_eFPGA_top.FrameData[123] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1244__I0 (.I(\Inst_eFPGA_top.FrameData[124] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1241__I1 (.I(\Inst_eFPGA_top.FrameData[124] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[28]  (.I(\Inst_eFPGA_top.FrameData[124] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1246__I0 (.I(\Inst_eFPGA_top.FrameData[125] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1244__I1 (.I(\Inst_eFPGA_top.FrameData[125] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[29]  (.I(\Inst_eFPGA_top.FrameData[125] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1248__I0 (.I(\Inst_eFPGA_top.FrameData[126] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1246__I1 (.I(\Inst_eFPGA_top.FrameData[126] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[30]  (.I(\Inst_eFPGA_top.FrameData[126] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1250__I0 (.I(\Inst_eFPGA_top.FrameData[127] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1248__I1 (.I(\Inst_eFPGA_top.FrameData[127] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[31]  (.I(\Inst_eFPGA_top.FrameData[127] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1034__I0 (.I(\Inst_eFPGA_top.FrameData[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1032__I1 (.I(\Inst_eFPGA_top.FrameData[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[1]  (.I(\Inst_eFPGA_top.FrameData[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1036__I0 (.I(\Inst_eFPGA_top.FrameData[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1034__I1 (.I(\Inst_eFPGA_top.FrameData[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[2]  (.I(\Inst_eFPGA_top.FrameData[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1038__I0 (.I(\Inst_eFPGA_top.FrameData[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1036__I1 (.I(\Inst_eFPGA_top.FrameData[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[3]  (.I(\Inst_eFPGA_top.FrameData[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1041__I0 (.I(\Inst_eFPGA_top.FrameData[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1038__I1 (.I(\Inst_eFPGA_top.FrameData[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[4]  (.I(\Inst_eFPGA_top.FrameData[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1047__I0 (.I(\Inst_eFPGA_top.FrameData[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1045__I1 (.I(\Inst_eFPGA_top.FrameData[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[7]  (.I(\Inst_eFPGA_top.FrameData[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1052__I0 (.I(\Inst_eFPGA_top.FrameData[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1050__I1 (.I(\Inst_eFPGA_top.FrameData[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[9]  (.I(\Inst_eFPGA_top.FrameData[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1054__I0 (.I(\Inst_eFPGA_top.FrameData[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1052__I1 (.I(\Inst_eFPGA_top.FrameData[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[10]  (.I(\Inst_eFPGA_top.FrameData[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1056__I0 (.I(\Inst_eFPGA_top.FrameData[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1054__I1 (.I(\Inst_eFPGA_top.FrameData[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[11]  (.I(\Inst_eFPGA_top.FrameData[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1059__I0 (.I(\Inst_eFPGA_top.FrameData[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1056__I1 (.I(\Inst_eFPGA_top.FrameData[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[12]  (.I(\Inst_eFPGA_top.FrameData[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1063__I0 (.I(\Inst_eFPGA_top.FrameData[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1061__I1 (.I(\Inst_eFPGA_top.FrameData[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[14]  (.I(\Inst_eFPGA_top.FrameData[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1065__I0 (.I(\Inst_eFPGA_top.FrameData[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1063__I1 (.I(\Inst_eFPGA_top.FrameData[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[15]  (.I(\Inst_eFPGA_top.FrameData[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1069__I0 (.I(\Inst_eFPGA_top.FrameData[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1065__I1 (.I(\Inst_eFPGA_top.FrameData[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[16]  (.I(\Inst_eFPGA_top.FrameData[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1071__I0 (.I(\Inst_eFPGA_top.FrameData[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1069__I1 (.I(\Inst_eFPGA_top.FrameData[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[17]  (.I(\Inst_eFPGA_top.FrameData[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1073__I0 (.I(\Inst_eFPGA_top.FrameData[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1071__I1 (.I(\Inst_eFPGA_top.FrameData[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[18]  (.I(\Inst_eFPGA_top.FrameData[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1075__I0 (.I(\Inst_eFPGA_top.FrameData[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1073__I1 (.I(\Inst_eFPGA_top.FrameData[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[19]  (.I(\Inst_eFPGA_top.FrameData[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1078__I0 (.I(\Inst_eFPGA_top.FrameData[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1075__I1 (.I(\Inst_eFPGA_top.FrameData[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[20]  (.I(\Inst_eFPGA_top.FrameData[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1080__I0 (.I(\Inst_eFPGA_top.FrameData[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1078__I1 (.I(\Inst_eFPGA_top.FrameData[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[21]  (.I(\Inst_eFPGA_top.FrameData[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1082__I0 (.I(\Inst_eFPGA_top.FrameData[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1080__I1 (.I(\Inst_eFPGA_top.FrameData[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[22]  (.I(\Inst_eFPGA_top.FrameData[54] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1096__I0 (.I(\Inst_eFPGA_top.FrameData[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1093__I1 (.I(\Inst_eFPGA_top.FrameData[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[28]  (.I(\Inst_eFPGA_top.FrameData[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1098__I0 (.I(\Inst_eFPGA_top.FrameData[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1096__I1 (.I(\Inst_eFPGA_top.FrameData[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[29]  (.I(\Inst_eFPGA_top.FrameData[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1100__I0 (.I(\Inst_eFPGA_top.FrameData[62] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1098__I1 (.I(\Inst_eFPGA_top.FrameData[62] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[30]  (.I(\Inst_eFPGA_top.FrameData[62] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1102__I0 (.I(\Inst_eFPGA_top.FrameData[63] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1100__I1 (.I(\Inst_eFPGA_top.FrameData[63] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_FrameData[31]  (.I(\Inst_eFPGA_top.FrameData[63] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1106__I0 (.I(\Inst_eFPGA_top.FrameData[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1102__I1 (.I(\Inst_eFPGA_top.FrameData[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[0]  (.I(\Inst_eFPGA_top.FrameData[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1108__I0 (.I(\Inst_eFPGA_top.FrameData[65] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1106__I1 (.I(\Inst_eFPGA_top.FrameData[65] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[1]  (.I(\Inst_eFPGA_top.FrameData[65] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1110__I0 (.I(\Inst_eFPGA_top.FrameData[66] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1108__I1 (.I(\Inst_eFPGA_top.FrameData[66] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[2]  (.I(\Inst_eFPGA_top.FrameData[66] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1115__I0 (.I(\Inst_eFPGA_top.FrameData[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1112__I1 (.I(\Inst_eFPGA_top.FrameData[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[4]  (.I(\Inst_eFPGA_top.FrameData[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1119__I0 (.I(\Inst_eFPGA_top.FrameData[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1117__I1 (.I(\Inst_eFPGA_top.FrameData[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[6]  (.I(\Inst_eFPGA_top.FrameData[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1121__I0 (.I(\Inst_eFPGA_top.FrameData[71] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1119__I1 (.I(\Inst_eFPGA_top.FrameData[71] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[7]  (.I(\Inst_eFPGA_top.FrameData[71] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1133__I0 (.I(\Inst_eFPGA_top.FrameData[76] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1130__I1 (.I(\Inst_eFPGA_top.FrameData[76] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[12]  (.I(\Inst_eFPGA_top.FrameData[76] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1135__I0 (.I(\Inst_eFPGA_top.FrameData[77] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1133__I1 (.I(\Inst_eFPGA_top.FrameData[77] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[13]  (.I(\Inst_eFPGA_top.FrameData[77] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1139__I0 (.I(\Inst_eFPGA_top.FrameData[79] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1137__I1 (.I(\Inst_eFPGA_top.FrameData[79] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[15]  (.I(\Inst_eFPGA_top.FrameData[79] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1161__I0 (.I(\Inst_eFPGA_top.FrameData[88] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1158__I1 (.I(\Inst_eFPGA_top.FrameData[88] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[24]  (.I(\Inst_eFPGA_top.FrameData[88] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1170__I0 (.I(\Inst_eFPGA_top.FrameData[92] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1167__I1 (.I(\Inst_eFPGA_top.FrameData[92] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[28]  (.I(\Inst_eFPGA_top.FrameData[92] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1172__I0 (.I(\Inst_eFPGA_top.FrameData[93] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1170__I1 (.I(\Inst_eFPGA_top.FrameData[93] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[29]  (.I(\Inst_eFPGA_top.FrameData[93] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1174__I0 (.I(\Inst_eFPGA_top.FrameData[94] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1172__I1 (.I(\Inst_eFPGA_top.FrameData[94] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[30]  (.I(\Inst_eFPGA_top.FrameData[94] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1176__I0 (.I(\Inst_eFPGA_top.FrameData[95] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1174__I1 (.I(\Inst_eFPGA_top.FrameData[95] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_FrameData[31]  (.I(\Inst_eFPGA_top.FrameData[95] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1180__I0 (.I(\Inst_eFPGA_top.FrameData[96] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1176__I1 (.I(\Inst_eFPGA_top.FrameData[96] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[0]  (.I(\Inst_eFPGA_top.FrameData[96] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1182__I0 (.I(\Inst_eFPGA_top.FrameData[97] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1180__I1 (.I(\Inst_eFPGA_top.FrameData[97] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[1]  (.I(\Inst_eFPGA_top.FrameData[97] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1184__I0 (.I(\Inst_eFPGA_top.FrameData[98] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1182__I1 (.I(\Inst_eFPGA_top.FrameData[98] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameData[2]  (.I(\Inst_eFPGA_top.FrameData[98] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[0]  (.I(\Inst_eFPGA_top.FrameSelect[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[10]  (.I(\Inst_eFPGA_top.FrameSelect[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[4]  (.I(\Inst_eFPGA_top.FrameSelect[112] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[5]  (.I(\Inst_eFPGA_top.FrameSelect[113] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[6]  (.I(\Inst_eFPGA_top.FrameSelect[114] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[7]  (.I(\Inst_eFPGA_top.FrameSelect[115] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[8]  (.I(\Inst_eFPGA_top.FrameSelect[116] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[9]  (.I(\Inst_eFPGA_top.FrameSelect[117] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[10]  (.I(\Inst_eFPGA_top.FrameSelect[118] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[11]  (.I(\Inst_eFPGA_top.FrameSelect[119] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[11]  (.I(\Inst_eFPGA_top.FrameSelect[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[12]  (.I(\Inst_eFPGA_top.FrameSelect[120] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[13]  (.I(\Inst_eFPGA_top.FrameSelect[121] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[14]  (.I(\Inst_eFPGA_top.FrameSelect[122] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[15]  (.I(\Inst_eFPGA_top.FrameSelect[123] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[16]  (.I(\Inst_eFPGA_top.FrameSelect[124] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[17]  (.I(\Inst_eFPGA_top.FrameSelect[125] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[18]  (.I(\Inst_eFPGA_top.FrameSelect[126] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[19]  (.I(\Inst_eFPGA_top.FrameSelect[127] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[12]  (.I(\Inst_eFPGA_top.FrameSelect[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[24]  (.I(\Inst_eFPGA_top.FrameSelect[132] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[25]  (.I(\Inst_eFPGA_top.FrameSelect[133] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[26]  (.I(\Inst_eFPGA_top.FrameSelect[134] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[27]  (.I(\Inst_eFPGA_top.FrameSelect[135] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[28]  (.I(\Inst_eFPGA_top.FrameSelect[136] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[29]  (.I(\Inst_eFPGA_top.FrameSelect[137] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[30]  (.I(\Inst_eFPGA_top.FrameSelect[138] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[31]  (.I(\Inst_eFPGA_top.FrameSelect[139] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[13]  (.I(\Inst_eFPGA_top.FrameSelect[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[32]  (.I(\Inst_eFPGA_top.FrameSelect[140] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[33]  (.I(\Inst_eFPGA_top.FrameSelect[141] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[34]  (.I(\Inst_eFPGA_top.FrameSelect[142] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_FrameStrobe[35]  (.I(\Inst_eFPGA_top.FrameSelect[143] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[0]  (.I(\Inst_eFPGA_top.FrameSelect[144] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[1]  (.I(\Inst_eFPGA_top.FrameSelect[145] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[14]  (.I(\Inst_eFPGA_top.FrameSelect[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[12]  (.I(\Inst_eFPGA_top.FrameSelect[156] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[14]  (.I(\Inst_eFPGA_top.FrameSelect[158] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[15]  (.I(\Inst_eFPGA_top.FrameSelect[159] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[15]  (.I(\Inst_eFPGA_top.FrameSelect[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[16]  (.I(\Inst_eFPGA_top.FrameSelect[160] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[17]  (.I(\Inst_eFPGA_top.FrameSelect[161] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[18]  (.I(\Inst_eFPGA_top.FrameSelect[162] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[19]  (.I(\Inst_eFPGA_top.FrameSelect[163] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[20]  (.I(\Inst_eFPGA_top.FrameSelect[164] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[21]  (.I(\Inst_eFPGA_top.FrameSelect[165] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[22]  (.I(\Inst_eFPGA_top.FrameSelect[166] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[23]  (.I(\Inst_eFPGA_top.FrameSelect[167] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[24]  (.I(\Inst_eFPGA_top.FrameSelect[168] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[25]  (.I(\Inst_eFPGA_top.FrameSelect[169] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[16]  (.I(\Inst_eFPGA_top.FrameSelect[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[26]  (.I(\Inst_eFPGA_top.FrameSelect[170] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[27]  (.I(\Inst_eFPGA_top.FrameSelect[171] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[28]  (.I(\Inst_eFPGA_top.FrameSelect[172] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[29]  (.I(\Inst_eFPGA_top.FrameSelect[173] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[30]  (.I(\Inst_eFPGA_top.FrameSelect[174] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[31]  (.I(\Inst_eFPGA_top.FrameSelect[175] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[32]  (.I(\Inst_eFPGA_top.FrameSelect[176] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[33]  (.I(\Inst_eFPGA_top.FrameSelect[177] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[34]  (.I(\Inst_eFPGA_top.FrameSelect[178] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_FrameStrobe[35]  (.I(\Inst_eFPGA_top.FrameSelect[179] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[17]  (.I(\Inst_eFPGA_top.FrameSelect[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[18]  (.I(\Inst_eFPGA_top.FrameSelect[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[19]  (.I(\Inst_eFPGA_top.FrameSelect[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[1]  (.I(\Inst_eFPGA_top.FrameSelect[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[20]  (.I(\Inst_eFPGA_top.FrameSelect[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[21]  (.I(\Inst_eFPGA_top.FrameSelect[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[22]  (.I(\Inst_eFPGA_top.FrameSelect[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[23]  (.I(\Inst_eFPGA_top.FrameSelect[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[24]  (.I(\Inst_eFPGA_top.FrameSelect[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[25]  (.I(\Inst_eFPGA_top.FrameSelect[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[26]  (.I(\Inst_eFPGA_top.FrameSelect[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[27]  (.I(\Inst_eFPGA_top.FrameSelect[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[28]  (.I(\Inst_eFPGA_top.FrameSelect[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[29]  (.I(\Inst_eFPGA_top.FrameSelect[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[2]  (.I(\Inst_eFPGA_top.FrameSelect[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[30]  (.I(\Inst_eFPGA_top.FrameSelect[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[31]  (.I(\Inst_eFPGA_top.FrameSelect[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[32]  (.I(\Inst_eFPGA_top.FrameSelect[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[33]  (.I(\Inst_eFPGA_top.FrameSelect[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[0]  (.I(\Inst_eFPGA_top.FrameSelect[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[1]  (.I(\Inst_eFPGA_top.FrameSelect[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[2]  (.I(\Inst_eFPGA_top.FrameSelect[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[3]  (.I(\Inst_eFPGA_top.FrameSelect[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[3]  (.I(\Inst_eFPGA_top.FrameSelect[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[4]  (.I(\Inst_eFPGA_top.FrameSelect[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[5]  (.I(\Inst_eFPGA_top.FrameSelect[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[6]  (.I(\Inst_eFPGA_top.FrameSelect[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[7]  (.I(\Inst_eFPGA_top.FrameSelect[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[8]  (.I(\Inst_eFPGA_top.FrameSelect[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[9]  (.I(\Inst_eFPGA_top.FrameSelect[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[10]  (.I(\Inst_eFPGA_top.FrameSelect[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[11]  (.I(\Inst_eFPGA_top.FrameSelect[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[4]  (.I(\Inst_eFPGA_top.FrameSelect[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[5]  (.I(\Inst_eFPGA_top.FrameSelect[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[28]  (.I(\Inst_eFPGA_top.FrameSelect[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[29]  (.I(\Inst_eFPGA_top.FrameSelect[65] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[30]  (.I(\Inst_eFPGA_top.FrameSelect[66] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[31]  (.I(\Inst_eFPGA_top.FrameSelect[67] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[32]  (.I(\Inst_eFPGA_top.FrameSelect[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[33]  (.I(\Inst_eFPGA_top.FrameSelect[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[6]  (.I(\Inst_eFPGA_top.FrameSelect[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[34]  (.I(\Inst_eFPGA_top.FrameSelect[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_FrameStrobe[35]  (.I(\Inst_eFPGA_top.FrameSelect[71] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[0]  (.I(\Inst_eFPGA_top.FrameSelect[72] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[1]  (.I(\Inst_eFPGA_top.FrameSelect[73] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[2]  (.I(\Inst_eFPGA_top.FrameSelect[74] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[3]  (.I(\Inst_eFPGA_top.FrameSelect[75] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[4]  (.I(\Inst_eFPGA_top.FrameSelect[76] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[5]  (.I(\Inst_eFPGA_top.FrameSelect[77] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[6]  (.I(\Inst_eFPGA_top.FrameSelect[78] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[7]  (.I(\Inst_eFPGA_top.FrameSelect[79] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[7]  (.I(\Inst_eFPGA_top.FrameSelect[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[12]  (.I(\Inst_eFPGA_top.FrameSelect[84] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[13]  (.I(\Inst_eFPGA_top.FrameSelect[85] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[14]  (.I(\Inst_eFPGA_top.FrameSelect[86] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[15]  (.I(\Inst_eFPGA_top.FrameSelect[87] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[16]  (.I(\Inst_eFPGA_top.FrameSelect[88] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[17]  (.I(\Inst_eFPGA_top.FrameSelect[89] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[8]  (.I(\Inst_eFPGA_top.FrameSelect[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[18]  (.I(\Inst_eFPGA_top.FrameSelect[90] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[19]  (.I(\Inst_eFPGA_top.FrameSelect[91] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[20]  (.I(\Inst_eFPGA_top.FrameSelect[92] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[21]  (.I(\Inst_eFPGA_top.FrameSelect[93] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[22]  (.I(\Inst_eFPGA_top.FrameSelect[94] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[23]  (.I(\Inst_eFPGA_top.FrameSelect[95] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[24]  (.I(\Inst_eFPGA_top.FrameSelect[96] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[25]  (.I(\Inst_eFPGA_top.FrameSelect[97] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[26]  (.I(\Inst_eFPGA_top.FrameSelect[98] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_FrameStrobe[27]  (.I(\Inst_eFPGA_top.FrameSelect[99] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_FrameStrobe[9]  (.I(\Inst_eFPGA_top.FrameSelect[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1532__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_A_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_B_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1528__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1516__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_A_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1527__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1515__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_B_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_A_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1511__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_B_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1518__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_A_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1529__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1517__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_B_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1526__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1514__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_A_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1513__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_B_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1522__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_A_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_I_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1509__I (.I(\Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_B_T_top ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[87].rs_and_A1  (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[88].rs_and_A1  (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[89].rs_and_A1  (.I(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[90].rs_and_A1  (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[91].rs_and_A1  (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[92].rs_and_A1  (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[93].rs_and_A1  (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[94].rs_and_A1  (.I(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[95].rs_and_A1  (.I(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[97].rs_and_A1  (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[112].rs_and_A1  (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[113].rs_and_A1  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[114].rs_and_A1  (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[115].rs_and_A1  (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[116].rs_and_A1  (.I(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[117].rs_and_A1  (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[118].rs_and_A1  (.I(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[119].rs_and_A1  (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[120].rs_and_A1  (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[122].rs_and_A1  (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[123].rs_and_A1  (.I(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[124].rs_and_A1  (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[125].rs_and_A1  (.I(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[126].rs_and_A1  (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[0].rs_and_A1  (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[127].rs_and_A1  (.I(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[132].rs_and_A1  (.I(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[133].rs_and_A1  (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[134].rs_and_A1  (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[135].rs_and_A1  (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[136].rs_and_A1  (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[1].rs_and_A1  (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[137].rs_and_A1  (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[138].rs_and_A1  (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[139].rs_and_A1  (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[140].rs_and_A1  (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[141].rs_and_A1  (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[142].rs_and_A1  (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[143].rs_and_A1  (.I(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[145].rs_and_A1  (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[2].rs_and_A1  (.I(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[148].rs_and_A1  (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[149].rs_and_A1  (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[150].rs_and_A1  (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[151].rs_and_A1  (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[152].rs_and_A1  (.I(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[153].rs_and_A1  (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[154].rs_and_A1  (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[155].rs_and_A1  (.I(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[156].rs_and_A1  (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[3].rs_and_A1  (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[157].rs_and_A1  (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[158].rs_and_A1  (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[159].rs_and_A1  (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[160].rs_and_A1  (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[161].rs_and_A1  (.I(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[163].rs_and_A1  (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[164].rs_and_A1  (.I(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[165].rs_and_A1  (.I(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[166].rs_and_A1  (.I(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[4].rs_and_A1  (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[167].rs_and_A1  (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[168].rs_and_A1  (.I(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[169].rs_and_A1  (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[170].rs_and_A1  (.I(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[171].rs_and_A1  (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[172].rs_and_A1  (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[173].rs_and_A1  (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[174].rs_and_A1  (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[175].rs_and_A1  (.I(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[176].rs_and_A1  (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[5].rs_and_A1  (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[177].rs_and_A1  (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[178].rs_and_A1  (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[179].rs_and_A1  (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[6].rs_and_A1  (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[7].rs_and_A1  (.I(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[8].rs_and_A1  (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[9].rs_and_A1  (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[10].rs_and_A1  (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[11].rs_and_A1  (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[12].rs_and_A1  (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[13].rs_and_A1  (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[14].rs_and_A1  (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[15].rs_and_A1  (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[16].rs_and_A1  (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[17].rs_and_A1  (.I(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[18].rs_and_A1  (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[19].rs_and_A1  (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[20].rs_and_A1  (.I(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[21].rs_and_A1  (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[22].rs_and_A1  (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[23].rs_and_A1  (.I(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[24].rs_and_A1  (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[25].rs_and_A1  (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[26].rs_and_A1  (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[27].rs_and_A1  (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[28].rs_and_A1  (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[29].rs_and_A1  (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[30].rs_and_A1  (.I(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[31].rs_and_A1  (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[32].rs_and_A1  (.I(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[33].rs_and_A1  (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[36].rs_and_A1  (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[37].rs_and_A1  (.I(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[38].rs_and_A1  (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[39].rs_and_A1  (.I(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[40].rs_and_A1  (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[42].rs_and_A1  (.I(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[44].rs_and_A1  (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[45].rs_and_A1  (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[65].rs_and_A1  (.I(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[67].rs_and_A1  (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[69].rs_and_A1  (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[70].rs_and_A1  (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[71].rs_and_A1  (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[72].rs_and_A1  (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[73].rs_and_A1  (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[74].rs_and_A1  (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[75].rs_and_A1  (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[76].rs_and_A1  (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[77].rs_and_A1  (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[78].rs_and_A1  (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[79].rs_and_A1  (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[86].rs_and_A1  (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1363__D (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1266__D (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1243__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1234__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1225__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1216__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1223__S (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1221__S (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1219__S (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1217__S (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1232__S (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1230__S (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1228__S (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1226__S (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1241__S (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1239__S (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1237__S (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1235__S (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1250__S (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1248__S (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1246__S (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1244__S (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1251__I (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0753__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0729__I (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0705__I (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0629__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1005__A4 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0989__A4 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0706__I (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0628__I (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0902__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0779__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0633__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0988__B (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0875__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0752__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0632__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0776__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0730__A3 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0708__A1 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0633__A2 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0690__I (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0676__I (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0661__I (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0634__I (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0660__A1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0656__A1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0651__A1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0645__A1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0977__B (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0677__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0663__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0637__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0658__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0654__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0649__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0643__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0970__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0969__B (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0648__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0642__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0969__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0967__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0966__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0642__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0657__A4 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0653__A4 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0648__A4 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0642__A4 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0693__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0678__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0664__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0643__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0874__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0775__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0644__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0756__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0732__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0710__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0645__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0972__A3 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0970__A3 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0653__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0647__I (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0696__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0681__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0667__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0649__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0879__I (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0782__I (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0650__I (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0757__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0733__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0711__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0651__A2 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0699__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0684__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0670__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0654__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0882__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0784__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0655__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0758__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0734__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0712__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0656__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0702__A1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0687__A1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0673__A1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0658__A2 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0884__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0786__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0659__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0759__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0735__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0713__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0660__A2 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0675__A1 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0672__A1 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0669__A1 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0666__A1 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0975__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0974__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0677__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0663__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0673__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0670__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0667__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0664__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0788__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0665__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0761__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0737__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0715__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0666__A2 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0792__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0668__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0762__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0738__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0716__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0669__A2 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0795__I (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0671__I (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0763__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0739__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0717__A1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0672__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0798__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0674__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0764__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0740__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0718__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0675__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0689__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0686__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0683__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0680__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0687__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0684__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0681__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0678__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0801__I (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0679__I (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0766__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0742__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0720__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0680__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0805__I (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0682__I (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0767__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0743__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0721__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0683__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0809__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0685__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0768__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0744__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0722__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0686__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0812__I (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0688__I (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0769__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0745__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0723__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0689__A2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0704__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0701__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0698__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0695__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0702__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0699__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0696__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0693__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0815__I (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0694__I (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0771__A1 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0747__A1 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0725__A1 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0695__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0819__I (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0697__I (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0772__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0748__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0726__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0698__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0822__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0700__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0773__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0749__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0727__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0701__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0825__I (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0703__I (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0774__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0750__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0728__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0704__A2 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0851__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0753__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0730__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0707__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0926__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0828__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0708__A2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0724__I (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0719__I (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0714__I (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0709__I (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0713__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0712__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0711__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0710__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0718__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0717__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0716__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0715__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0723__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0722__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0721__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0720__A2 (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0983__B (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0949__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0851__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0730__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0746__I (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0741__I (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0736__I (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0731__I (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0735__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0734__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0733__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0732__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0740__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0739__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0738__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0737__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0750__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0749__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0748__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0747__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0986__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0875__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0752__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0851__A3 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0828__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0779__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0754__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0876__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0776__A2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0754__A2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0770__I (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0765__I (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0760__I (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0755__I (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0759__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0758__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0757__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0756__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0764__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0763__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0762__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0761__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0853__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0830__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0781__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0778__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0956__I (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0924__I (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0862__I (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0777__I (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0848__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0834__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0808__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0778__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0817__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0803__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0790__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0780__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0787__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0785__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0783__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0781__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0854__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0831__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0808__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0783__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0855__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0834__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0832__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0785__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0856__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0848__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0833__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0787__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0933__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0909__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0887__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0789__I (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0863__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0858__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0836__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0791__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0800__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0797__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0794__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0791__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0934__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0910__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0888__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0793__I (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0881__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0859__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0837__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0794__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0935__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0912__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0896__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0796__I (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0889__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0860__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0838__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0797__A1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0936__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0913__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0911__A1 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0799__I (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0890__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0861__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0839__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0800__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0938__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0925__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0915__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0802__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0892__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0865__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0841__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0804__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0814__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0811__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0807__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0804__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0940__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0939__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0916__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0806__I (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0893__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0866__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0842__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0807__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0954__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0941__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0917__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0810__I (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0894__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0867__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0843__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0811__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0955__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0942__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0918__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0813__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0895__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0868__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0844__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0814__A1 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0957__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0944__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0920__A1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0816__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0898__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0870__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0846__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0818__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0827__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0824__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0821__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0818__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0958__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0945__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0921__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0820__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0899__A1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0871__A1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0847__A1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0821__A1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0959__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0946__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0922__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0823__I (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0900__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0872__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0849__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0824__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0960__A1 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0947__A1 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0923__A1 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0826__I (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0901__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0873__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0850__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0827__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0845__I (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0840__I (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0835__I (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0829__I (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0833__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0832__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0831__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0830__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0839__A2 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0838__A2 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0837__A2 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0836__A2 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0844__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0843__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0842__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0841__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0850__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0849__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0847__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0846__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0869__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0864__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0857__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0852__I (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0856__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0855__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0854__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0853__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0861__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0860__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0859__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0858__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0911__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0896__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0881__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0863__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0868__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0867__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0866__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0865__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0873__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0872__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0871__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0870__A2 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0950__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0928__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0904__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0878__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0949__A3 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0926__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0902__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0876__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0897__I (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0891__I (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0886__I (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0877__I (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0885__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0883__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0880__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0878__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0951__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0929__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0905__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0880__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0952__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0930__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0906__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0883__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0953__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0931__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0907__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0885__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0895__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0894__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0893__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0892__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0901__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0900__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0899__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0898__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0919__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0914__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0908__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0903__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0907__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0906__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0905__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0904__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0913__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0912__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0910__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0909__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0918__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0917__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0916__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0915__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0923__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0922__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0921__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0920__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0955__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0954__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0940__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0925__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0943__I (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0937__I (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0932__I (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0927__I (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0931__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0930__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0929__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0928__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0936__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0935__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0934__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0933__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0942__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0941__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0939__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0938__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0947__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0946__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0945__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0944__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0983__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0982__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0981__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0949__A2 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0953__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0952__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0951__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0950__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0960__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0959__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0958__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0957__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1016__B (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1002__B (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0998__B (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0965__I (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1027__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0981__B (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0974__B (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0966__B (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1013__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0994__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0987__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0971__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1011__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1007__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0977__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0971__A3 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0990__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0984__A4 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0973__I (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1009__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0991__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0985__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0980__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0997__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0990__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0984__A3 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0979__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0983__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0982__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0981__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0980__A3 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0997__A3 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0990__A3 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0999__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0993__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0991__A3 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1006__A4 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0998__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0996__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0993__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1006__A3 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0999__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0998__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0996__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1004__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1003__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1002__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1000__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1006__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1004__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1003__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1002__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1021__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1016__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1015__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1012__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1025__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1022__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1012__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1023__A2 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1025__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1022__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1023__A3 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1141__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1104__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1067__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1030__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1058__I (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1049__I (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1040__I (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1031__I (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1056__S (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1054__S (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1052__S (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1050__S (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1065__S (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1063__S (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1061__S (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1059__S (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1095__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1086__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1077__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1068__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1084__S (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1082__S (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1080__S (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1078__S (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1093__S (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1091__S (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1089__S (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1087__S (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1102__S (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1100__S (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1098__S (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1096__S (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1132__I (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1123__I (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1114__I (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1105__I (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1112__S (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1110__S (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1108__S (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1106__S (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1121__S (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1119__S (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1117__S (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1115__S (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1130__S (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1128__S (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1126__S (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1124__S (.I(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1169__I (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1160__I (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1151__I (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1142__I (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1149__S (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1147__S (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1145__S (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1143__S (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1176__S (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1174__S (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1172__S (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1170__S (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1206__I (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1197__I (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1188__I (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1179__I (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1186__S (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1184__S (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1182__S (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1180__S (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1195__S (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1193__S (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1191__S (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1189__S (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1204__S (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1202__S (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1200__S (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1198__S (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1213__S (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1211__S (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1209__S (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1207__S (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1006__A1 (.I(\fstb_ctr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1004__B (.I(\fstb_ctr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0640__A3 (.I(\fstb_ctr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0972__A2 (.I(\fstb_ctr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0652__I (.I(\fstb_ctr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0638__I (.I(\fstb_ctr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1005__A3 (.I(\fstb_ctr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0989__A3 (.I(\fstb_ctr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0626__I (.I(\fstb_ctr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1005__A1 (.I(\fstb_ctr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0989__A1 (.I(\fstb_ctr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0630__I (.I(\fstb_ctr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(io_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_in[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(io_in[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(io_in[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_0_io_in[5]_I  (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_2_3_0_io_in[5]_I  (.I(clknet_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_2_2_0_io_in[5]_I  (.I(clknet_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_2_1_0_io_in[5]_I  (.I(clknet_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_2_0_0_io_in[5]_I  (.I(clknet_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(la_data_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(la_data_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[9].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[99].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[98].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[97].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[96].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[95].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[94].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[93].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[92].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[91].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[90].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[8].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[89].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[88].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[87].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[86].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[85].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[84].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[83].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[82].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[81].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[80].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[7].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[79].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[78].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[77].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[76].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[75].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[74].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[73].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[72].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[71].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[70].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[6].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[69].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[68].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[67].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[66].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[65].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[64].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[63].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[62].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[61].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[60].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[5].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[59].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[58].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[57].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[56].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[55].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[54].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[53].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[52].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[51].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[50].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[4].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[49].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[48].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[47].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[46].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[45].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[44].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[43].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[42].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[41].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[40].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[3].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[39].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[38].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[37].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[36].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[35].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[34].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[33].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[32].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[31].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[30].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[2].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[29].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[28].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[27].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[26].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[25].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[24].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[23].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[22].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[21].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[20].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[1].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[19].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[18].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[17].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[179].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[178].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[177].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[176].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[175].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[174].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[173].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[172].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[171].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[170].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[16].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[169].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[168].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[167].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[166].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[165].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[164].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[163].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[162].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[161].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[160].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[15].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[159].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[158].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[157].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[156].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[155].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[154].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[153].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[152].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[151].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[150].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[14].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[149].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[148].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[147].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[146].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[145].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[144].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[143].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[142].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[141].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[140].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[13].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[139].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[138].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[137].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[136].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[135].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[134].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[133].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[132].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[131].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[130].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[12].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[129].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[128].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[127].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[126].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[125].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[124].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[123].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[122].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[121].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[120].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[11].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[119].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[118].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[117].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[116].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[115].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[114].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[113].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[112].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[111].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[110].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[10].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[109].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[108].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[107].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[106].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[105].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[104].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[103].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[102].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[101].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[100].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_frame_ands[0].rs_and_A2  (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_UserCLK  (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_sram_test1_i_WL (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_sram_test0_i_WL (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_sram_test0_i_BLP (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0961__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_sram_test1_i_BLP (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0962__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_B_O_top  (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y3_E_IO_A_O_top  (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_B_O_top  (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_A_O_top  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_E_IO_B_O_top  (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y2_E_IO_A_O_top  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_B_O_top  (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y2_W_IO_A_O_top  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_E_IO_B_O_top  (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X4Y1_E_IO_A_O_top  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_B_O_top  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y1_W_IO_A_O_top  (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1215__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1178__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1029__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1250__I1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1023__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0976__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0968__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0964__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0972__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0963__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_sram_test0_i_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_sram_test1_i_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output46_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output47_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output48_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_sram_test0_i_O (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_sram_test1_i_O (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X3Y4_S_term_single_OutputEnable  (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_OutputEnable  (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_OutputEnable  (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X0Y3_W_IO_UserCLK  (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_1_0_io_in[5]_I  (.I(clknet_2_0_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_0_0_io_in[5]_I  (.I(clknet_2_0_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_3_0_io_in[5]_I  (.I(clknet_2_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_2_0_io_in[5]_I  (.I(clknet_2_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_5_0_io_in[5]_I  (.I(clknet_2_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_4_0_io_in[5]_I  (.I(clknet_2_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_7_0_io_in[5]_I  (.I(clknet_2_3_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_6_0_io_in[5]_I  (.I(clknet_2_3_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_1_0_io_in[5]_I  (.I(clknet_3_0_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_0_0_io_in[5]_I  (.I(clknet_3_0_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_3_0_io_in[5]_I  (.I(clknet_3_1_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_2_0_io_in[5]_I  (.I(clknet_3_1_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_4_1_io_in[5]_I  (.I(clknet_3_4_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_9_0_io_in[5]_I  (.I(clknet_3_4_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_8_0_io_in[5]_I  (.I(clknet_3_4_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_5_1_io_in[5]_I  (.I(clknet_3_5_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_11_0_io_in[5]_I  (.I(clknet_3_5_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_10_0_io_in[5]_I  (.I(clknet_3_5_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_13_0_io_in[5]_I  (.I(clknet_3_6_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_12_0_io_in[5]_I  (.I(clknet_3_6_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_15_0_io_in[5]_I  (.I(clknet_3_7_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_4_14_0_io_in[5]_I  (.I(clknet_3_7_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1333__CLK (.I(clknet_4_0_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1334__CLK (.I(clknet_4_0_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1335__CLK (.I(clknet_4_0_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1336__CLK (.I(clknet_4_0_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1337__CLK (.I(clknet_4_0_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1338__CLK (.I(clknet_4_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1339__CLK (.I(clknet_4_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1340__CLK (.I(clknet_4_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1341__CLK (.I(clknet_4_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1342__CLK (.I(clknet_4_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1343__CLK (.I(clknet_4_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1345__CLK (.I(clknet_4_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1350__CLK (.I(clknet_4_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1351__CLK (.I(clknet_4_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1352__CLK (.I(clknet_4_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1353__CLK (.I(clknet_4_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1354__CLK (.I(clknet_4_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1355__CLK (.I(clknet_4_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1356__CLK (.I(clknet_4_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1357__CLK (.I(clknet_4_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1358__CLK (.I(clknet_4_2_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1332__CLK (.I(clknet_4_3_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1344__CLK (.I(clknet_4_3_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1346__CLK (.I(clknet_4_3_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1347__CLK (.I(clknet_4_3_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1348__CLK (.I(clknet_4_3_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1349__CLK (.I(clknet_4_3_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X1Y4_S_term_single_UserCLK  (.I(clknet_4_4_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1257__CLK (.I(clknet_4_4_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1258__CLK (.I(clknet_4_4_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1267__CLK (.I(clknet_4_4_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1252__CLK (.I(clknet_4_5_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1254__CLK (.I(clknet_4_5_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1259__CLK (.I(clknet_4_5_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1261__CLK (.I(clknet_4_5_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_Inst_eFPGA_top.Inst_eFPGA.Tile_X2Y4_S_term_single_UserCLK  (.I(clknet_4_6_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1253__CLK (.I(clknet_4_6_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1260__CLK (.I(clknet_4_6_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1263__CLK (.I(clknet_4_6_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1265__CLK (.I(clknet_4_6_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_opt_1_0_io_in[5]_I  (.I(clknet_4_7_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1255__CLK (.I(clknet_4_7_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1256__CLK (.I(clknet_4_7_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1262__CLK (.I(clknet_4_7_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1264__CLK (.I(clknet_4_7_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1266__CLK (.I(clknet_4_7_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1277__CLK (.I(clknet_4_8_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1278__CLK (.I(clknet_4_8_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1279__CLK (.I(clknet_4_8_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1280__CLK (.I(clknet_4_8_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1282__CLK (.I(clknet_4_8_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1286__CLK (.I(clknet_4_8_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1299__CLK (.I(clknet_4_8_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1324__CLK (.I(clknet_4_9_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1325__CLK (.I(clknet_4_9_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1326__CLK (.I(clknet_4_9_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1327__CLK (.I(clknet_4_9_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1329__CLK (.I(clknet_4_9_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1268__CLK (.I(clknet_4_10_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1269__CLK (.I(clknet_4_10_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1272__CLK (.I(clknet_4_10_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1275__CLK (.I(clknet_4_10_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1281__CLK (.I(clknet_4_10_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1283__CLK (.I(clknet_4_10_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1284__CLK (.I(clknet_4_10_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1273__CLK (.I(clknet_4_11_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1287__CLK (.I(clknet_4_11_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1289__CLK (.I(clknet_4_11_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1290__CLK (.I(clknet_4_11_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1291__CLK (.I(clknet_4_11_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1292__CLK (.I(clknet_4_11_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1293__CLK (.I(clknet_4_11_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1294__CLK (.I(clknet_4_11_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1298__CLK (.I(clknet_4_11_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1300__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1306__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1307__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1308__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1309__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1310__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1311__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1312__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1313__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1314__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1315__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1316__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1317__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1318__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1331__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1363__CLK (.I(clknet_4_12_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1301__CLK (.I(clknet_4_13_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1302__CLK (.I(clknet_4_13_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1303__CLK (.I(clknet_4_13_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1304__CLK (.I(clknet_4_13_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1305__CLK (.I(clknet_4_13_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1359__CLK (.I(clknet_4_13_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1360__CLK (.I(clknet_4_13_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1361__CLK (.I(clknet_4_13_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1362__CLK (.I(clknet_4_13_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1270__CLK (.I(clknet_4_14_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1271__CLK (.I(clknet_4_14_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1274__CLK (.I(clknet_4_14_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1276__CLK (.I(clknet_4_14_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1285__CLK (.I(clknet_4_14_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1288__CLK (.I(clknet_4_14_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1295__CLK (.I(clknet_4_14_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1296__CLK (.I(clknet_4_14_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1297__CLK (.I(clknet_4_14_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1319__CLK (.I(clknet_4_15_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1320__CLK (.I(clknet_4_15_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1321__CLK (.I(clknet_4_15_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1322__CLK (.I(clknet_4_15_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1323__CLK (.I(clknet_4_15_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1328__CLK (.I(clknet_4_15_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1330__CLK (.I(clknet_4_15_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_opt_1_1_io_in[5]_I  (.I(clknet_opt_1_0_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_opt_1_2_io_in[5]_I  (.I(clknet_opt_1_1_io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_247_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_248_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_249_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_250_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_251_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_252_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_253_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_254_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_254_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_260_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_262_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_262_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_263_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_268_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_268_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_269_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_269_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_270_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_270_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_271_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_272_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_273_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_274_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_274_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_274_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_275_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_278_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_279_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_280_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_281_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_282_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_282_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_283_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_284_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_288_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_289_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_290_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_291_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_292_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_293_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_293_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_294_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_294_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_295_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_295_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_296_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_297_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_297_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_298_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_299_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_300_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_301_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_301_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_302_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_303_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_303_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_304_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_305_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_305_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_306_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_307_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_307_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_308_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_309_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_309_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_310_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_311_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_311_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_312_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_314_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_314_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_315_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_316_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_316_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_318_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_319_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_319_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_320_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_320_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_321_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_322_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_323_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_323_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_325_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_326_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_328_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_328_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_329_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_329_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_330_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_330_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_330_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_330_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_331_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_331_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_331_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_331_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_331_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_331_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_332_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_332_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_333_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_333_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_333_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_333_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_333_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_333_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_333_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_334_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_334_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_334_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_335_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_335_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_336_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_337_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_337_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_337_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_337_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_337_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_338_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_338_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_338_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_338_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_338_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_338_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_339_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_339_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_339_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_339_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_339_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_340_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_341_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_341_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_342_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_342_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_342_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_342_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_342_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_342_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_343_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_343_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_343_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_344_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_345_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_345_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_345_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_346_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_346_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_346_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_346_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_346_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_346_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_346_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_346_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_346_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_346_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_347_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_347_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_348_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_348_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_348_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_348_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_348_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_348_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_348_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_348_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_348_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_349_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_349_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_349_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_350_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_350_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_351_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_351_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_351_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_351_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_351_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_351_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_351_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_352_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_352_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_352_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_352_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_352_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_352_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_353_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_353_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_353_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_353_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_353_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_353_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_354_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_354_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_354_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_355_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_355_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_355_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_355_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_355_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_355_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_355_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_356_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_356_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_356_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_356_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_356_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_356_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_356_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_356_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_357_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_357_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_357_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_357_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_357_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_358_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_358_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_358_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_358_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_358_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_358_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_358_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_359_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_359_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_359_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_360_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_360_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_360_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_361_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_361_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_361_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_361_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_362_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_362_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_362_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_362_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_362_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_362_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_363_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_363_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_363_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_363_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_363_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_363_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_363_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_363_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_364_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_364_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_364_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_365_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_365_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_365_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_365_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_366_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_366_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_366_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_367_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_367_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_367_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_368_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_368_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_369_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_369_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_369_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_370_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_370_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_370_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_371_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_371_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_371_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_372_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_372_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_373_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_374_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_374_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_374_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_374_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_374_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_374_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_374_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_375_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_375_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_376_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_376_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_376_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_376_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_376_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_376_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_376_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_377_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_377_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_377_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_378_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_378_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_378_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_378_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_378_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_378_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_378_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_379_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_379_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_380_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_380_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_380_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_380_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_380_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_380_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_380_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_381_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_381_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_382_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_382_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_382_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_382_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_382_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_382_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_382_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_383_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_383_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_384_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_384_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_384_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_384_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_384_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_384_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_384_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_385_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_385_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_386_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_386_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_386_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_386_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_386_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_386_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_386_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_387_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_387_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_388_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_388_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_388_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_388_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_388_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_388_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_388_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_389_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_389_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_390_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_390_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_390_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_390_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_390_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_390_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_390_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_391_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_391_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_392_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_392_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_392_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_392_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_392_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_392_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_392_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_393_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_393_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_394_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_394_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_394_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_394_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_394_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_394_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_394_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_395_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_395_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_396_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_396_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_396_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_396_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_396_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_396_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_396_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_397_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_397_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_398_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_398_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_398_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_398_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_398_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_398_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_398_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_399_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_399_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_400_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_400_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_400_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_400_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_400_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_400_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_400_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_401_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_401_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_402_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_402_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_402_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_402_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_402_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_402_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_402_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_403_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_403_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_404_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_404_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_404_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_404_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_404_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_404_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_404_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_405_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_405_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_406_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_406_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_406_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_406_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_406_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_406_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_406_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_407_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_407_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_408_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_408_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_408_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_408_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_408_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_408_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_408_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_409_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_409_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_410_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_410_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_410_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_410_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_410_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_410_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_410_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_411_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_411_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_412_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_412_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_412_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_412_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_412_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_412_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_412_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_413_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_413_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_414_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_414_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_414_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_414_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_414_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_414_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_414_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_415_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_415_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_416_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_416_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_416_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_416_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_416_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_416_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_416_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_417_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_417_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_418_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_418_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_418_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_418_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_418_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_418_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_418_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_419_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_419_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_420_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_420_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_420_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_420_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_420_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_420_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_421_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_421_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_421_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_421_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_421_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_421_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_421_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_422_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_422_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_422_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_422_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_422_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_422_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_423_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_423_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_423_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_423_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_423_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_423_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_423_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_423_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_423_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_423_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_423_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_423_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_3008 ();
 assign io_oeb[0] = net185;
 assign io_oeb[10] = net195;
 assign io_oeb[11] = net51;
 assign io_oeb[12] = net52;
 assign io_oeb[13] = net53;
 assign io_oeb[14] = net54;
 assign io_oeb[15] = net55;
 assign io_oeb[16] = net56;
 assign io_oeb[17] = net57;
 assign io_oeb[18] = net58;
 assign io_oeb[19] = net59;
 assign io_oeb[1] = net186;
 assign io_oeb[20] = net60;
 assign io_oeb[21] = net61;
 assign io_oeb[22] = net62;
 assign io_oeb[23] = net63;
 assign io_oeb[24] = net64;
 assign io_oeb[25] = net65;
 assign io_oeb[2] = net187;
 assign io_oeb[3] = net188;
 assign io_oeb[4] = net189;
 assign io_oeb[5] = net190;
 assign io_oeb[6] = net191;
 assign io_oeb[7] = net192;
 assign io_oeb[8] = net193;
 assign io_oeb[9] = net194;
 assign io_out[0] = net66;
 assign io_out[10] = net76;
 assign io_out[11] = net77;
 assign io_out[14] = net78;
 assign io_out[15] = net79;
 assign io_out[16] = net80;
 assign io_out[17] = net81;
 assign io_out[18] = net82;
 assign io_out[19] = net83;
 assign io_out[1] = net67;
 assign io_out[20] = net84;
 assign io_out[21] = net85;
 assign io_out[22] = net86;
 assign io_out[23] = net87;
 assign io_out[24] = net88;
 assign io_out[25] = net89;
 assign io_out[2] = net68;
 assign io_out[3] = net69;
 assign io_out[4] = net70;
 assign io_out[5] = net71;
 assign io_out[6] = net72;
 assign io_out[7] = net73;
 assign io_out[8] = net74;
 assign io_out[9] = net75;
 assign la_data_out[10] = net98;
 assign la_data_out[11] = net99;
 assign la_data_out[12] = net100;
 assign la_data_out[13] = net101;
 assign la_data_out[14] = net102;
 assign la_data_out[15] = net103;
 assign la_data_out[16] = net104;
 assign la_data_out[17] = net105;
 assign la_data_out[18] = net106;
 assign la_data_out[19] = net107;
 assign la_data_out[20] = net108;
 assign la_data_out[21] = net109;
 assign la_data_out[22] = net110;
 assign la_data_out[23] = net111;
 assign la_data_out[24] = net112;
 assign la_data_out[25] = net113;
 assign la_data_out[26] = net114;
 assign la_data_out[27] = net115;
 assign la_data_out[28] = net116;
 assign la_data_out[29] = net117;
 assign la_data_out[2] = net90;
 assign la_data_out[30] = net118;
 assign la_data_out[31] = net119;
 assign la_data_out[32] = net120;
 assign la_data_out[33] = net121;
 assign la_data_out[34] = net122;
 assign la_data_out[35] = net123;
 assign la_data_out[36] = net124;
 assign la_data_out[37] = net125;
 assign la_data_out[38] = net126;
 assign la_data_out[39] = net127;
 assign la_data_out[3] = net91;
 assign la_data_out[40] = net128;
 assign la_data_out[41] = net129;
 assign la_data_out[42] = net130;
 assign la_data_out[43] = net131;
 assign la_data_out[44] = net132;
 assign la_data_out[45] = net133;
 assign la_data_out[46] = net134;
 assign la_data_out[47] = net135;
 assign la_data_out[48] = net136;
 assign la_data_out[49] = net137;
 assign la_data_out[4] = net92;
 assign la_data_out[50] = net138;
 assign la_data_out[51] = net139;
 assign la_data_out[52] = net140;
 assign la_data_out[53] = net141;
 assign la_data_out[54] = net142;
 assign la_data_out[55] = net143;
 assign la_data_out[56] = net144;
 assign la_data_out[57] = net145;
 assign la_data_out[58] = net146;
 assign la_data_out[59] = net147;
 assign la_data_out[5] = net93;
 assign la_data_out[60] = net148;
 assign la_data_out[61] = net149;
 assign la_data_out[62] = net150;
 assign la_data_out[63] = net151;
 assign la_data_out[6] = net94;
 assign la_data_out[7] = net95;
 assign la_data_out[8] = net96;
 assign la_data_out[9] = net97;
 assign wbs_ack_o = net152;
 assign wbs_dat_o[0] = net153;
 assign wbs_dat_o[10] = net163;
 assign wbs_dat_o[11] = net164;
 assign wbs_dat_o[12] = net165;
 assign wbs_dat_o[13] = net166;
 assign wbs_dat_o[14] = net167;
 assign wbs_dat_o[15] = net168;
 assign wbs_dat_o[16] = net169;
 assign wbs_dat_o[17] = net170;
 assign wbs_dat_o[18] = net171;
 assign wbs_dat_o[19] = net172;
 assign wbs_dat_o[1] = net154;
 assign wbs_dat_o[20] = net173;
 assign wbs_dat_o[21] = net174;
 assign wbs_dat_o[22] = net175;
 assign wbs_dat_o[23] = net176;
 assign wbs_dat_o[24] = net177;
 assign wbs_dat_o[25] = net178;
 assign wbs_dat_o[26] = net179;
 assign wbs_dat_o[27] = net180;
 assign wbs_dat_o[28] = net181;
 assign wbs_dat_o[29] = net182;
 assign wbs_dat_o[2] = net155;
 assign wbs_dat_o[30] = net183;
 assign wbs_dat_o[31] = net184;
 assign wbs_dat_o[3] = net156;
 assign wbs_dat_o[4] = net157;
 assign wbs_dat_o[5] = net158;
 assign wbs_dat_o[6] = net159;
 assign wbs_dat_o[7] = net160;
 assign wbs_dat_o[8] = net161;
 assign wbs_dat_o[9] = net162;
endmodule

